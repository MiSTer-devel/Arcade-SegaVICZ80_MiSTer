// The following code is a copy of the T48 core by Arnim Läuger which has been automatically converted to Verilog for ease of simulation
// https://github.com/devsaurus/t48

`timescale 1ps / 1ps

module t48_decoder_1
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  ea_i,
   input  ale_i,
   input  int_n_i,
   input  [7:0] data_i,
   input  alu_carry_i,
   input  alu_da_overflow_i,
   input  [2:0] clk_mstate_i,
   input  clk_second_cycle_i,
   input  cnd_take_branch_i,
   input  psw_carry_i,
   input  psw_aux_carry_i,
   input  psw_f0_i,
   input  tim_overflow_i,
   output t0_dir_o,
   output [7:0] data_o,
   output alu_write_accu_o,
   output alu_write_shadow_o,
   output alu_write_temp_reg_o,
   output alu_read_alu_o,
   output bus_write_bus_o,
   output bus_read_bus_o,
   output dm_write_dmem_addr_o,
   output dm_write_dmem_o,
   output dm_read_dmem_o,
   output p1_write_p1_o,
   output p1_read_p1_o,
   output p2_write_p2_o,
   output p2_write_exp_o,
   output p2_read_p2_o,
   output p2_read_exp_o,
   output pm_write_pcl_o,
   output pm_read_pcl_o,
   output pm_write_pch_o,
   output pm_read_pch_o,
   output pm_read_pmem_o,
   output psw_read_psw_o,
   output psw_read_sp_o,
   output psw_write_psw_o,
   output psw_write_sp_o,
   output [3:0] alu_op_o,
   output alu_use_carry_o,
   output alu_da_high_o,
   output alu_accu_low_o,
   output alu_p06_temp_reg_o,
   output alu_p60_temp_reg_o,
   output bus_output_pcl_o,
   output bus_bidir_bus_o,
   output clk_multi_cycle_o,
   output clk_assert_psen_o,
   output clk_assert_prog_o,
   output clk_assert_rd_o,
   output clk_assert_wr_o,
   output cnd_compute_take_o,
   output [3:0] cnd_branch_cond_o,
   output [2:0] cnd_comp_value_o,
   output cnd_f1_o,
   output cnd_tf_o,
   output [1:0] dm_addr_type_o,
   output p1_read_reg_o,
   output p2_read_reg_o,
   output p2_output_pch_o,
   output pm_inc_pc_o,
   output pm_write_pmem_addr_o,
   output [1:0] pm_addr_type_o,
   output psw_special_data_o,
   output psw_inc_stackp_o,
   output psw_dec_stackp_o,
   output psw_write_carry_o,
   output psw_write_aux_carry_o,
   output psw_write_f0_o,
   output psw_write_bs_o,
   output tim_read_timer_o,
   output tim_write_timer_o,
   output tim_start_t_o,
   output tim_start_cnt_o,
   output tim_stop_tcnt_o);
  wire opc_multi_cycle_s;
  wire opc_read_bus_s;
  wire opc_inj_int_s;
  wire [7:0] opc_opcode_q;
  wire [5:0] opc_mnemonic_s;
  wire last_cycle_s;
  wire assert_psen_s;
  wire branch_taken_s;
  wire branch_taken_q;
  wire pm_inc_pc_s;
  wire pm_write_pmem_addr_s;
  wire add_inc_pc_s;
  wire add_write_pmem_addr_s;
  wire clear_f1_s;
  wire cpl_f1_s;
  wire f1_q;
  wire clear_mb_s;
  wire set_mb_s;
  wire mb_q;
  wire ent0_clk_s;
  wire t0_dir_q;
  wire [7:0] data_s;
  wire read_dec_s;
  wire tf_s;
  wire bus_read_bus_s;
  wire add_read_bus_s;
  wire dm_write_dmem_s;
  wire p2_output_exp_s;
  wire movx_first_cycle_s;
  wire jtf_executed_s;
  wire en_tcnti_s;
  wire dis_tcnti_s;
  wire en_i_s;
  wire dis_i_s;
  wire tim_int_s;
  wire retr_executed_s;
  wire int_executed_s;
  wire int_pending_s;
  wire int_in_progress_s;
  wire [6:0] mnemonic_rec_s;
  wire [5:0] mnemonic_q;
  wire n1179_o;
  wire n1181_o;
  wire n1182_o;
  wire n1184_o;
  wire n1185_o;
  wire n1187_o;
  wire n1188_o;
  wire n1190_o;
  wire n1191_o;
  wire n1193_o;
  wire n1194_o;
  wire n1196_o;
  wire n1197_o;
  wire n1199_o;
  wire n1200_o;
  wire n1202_o;
  wire n1203_o;
  wire n1205_o;
  wire n1206_o;
  wire n1208_o;
  wire n1209_o;
  wire n1211_o;
  wire n1212_o;
  wire n1214_o;
  wire n1215_o;
  wire n1217_o;
  wire n1218_o;
  wire n1220_o;
  wire n1221_o;
  wire n1223_o;
  wire n1224_o;
  wire n1226_o;
  wire n1227_o;
  wire n1229_o;
  wire n1230_o;
  wire n1232_o;
  wire n1233_o;
  wire n1235_o;
  wire n1236_o;
  wire n1238_o;
  wire n1240_o;
  wire n1241_o;
  wire n1243_o;
  wire n1245_o;
  wire n1246_o;
  wire n1248_o;
  wire n1249_o;
  wire n1251_o;
  wire n1252_o;
  wire n1254_o;
  wire n1255_o;
  wire n1257_o;
  wire n1258_o;
  wire n1260_o;
  wire n1261_o;
  wire n1263_o;
  wire n1264_o;
  wire n1266_o;
  wire n1267_o;
  wire n1269_o;
  wire n1270_o;
  wire n1272_o;
  wire n1274_o;
  wire n1276_o;
  wire n1277_o;
  wire n1279_o;
  wire n1280_o;
  wire n1282_o;
  wire n1284_o;
  wire n1285_o;
  wire n1287_o;
  wire n1288_o;
  wire n1290_o;
  wire n1291_o;
  wire n1293_o;
  wire n1294_o;
  wire n1296_o;
  wire n1297_o;
  wire n1299_o;
  wire n1300_o;
  wire n1302_o;
  wire n1303_o;
  wire n1305_o;
  wire n1307_o;
  wire n1309_o;
  wire n1311_o;
  wire n1312_o;
  wire n1314_o;
  wire n1316_o;
  wire n1318_o;
  wire n1320_o;
  wire n1321_o;
  wire n1323_o;
  wire n1325_o;
  wire n1327_o;
  wire n1328_o;
  wire n1330_o;
  wire n1331_o;
  wire n1333_o;
  wire n1334_o;
  wire n1336_o;
  wire n1337_o;
  wire n1339_o;
  wire n1340_o;
  wire n1342_o;
  wire n1343_o;
  wire n1345_o;
  wire n1346_o;
  wire n1348_o;
  wire n1349_o;
  wire n1351_o;
  wire n1353_o;
  wire n1354_o;
  wire n1356_o;
  wire n1358_o;
  wire n1359_o;
  wire n1361_o;
  wire n1363_o;
  wire n1364_o;
  wire n1366_o;
  wire n1367_o;
  wire n1369_o;
  wire n1370_o;
  wire n1372_o;
  wire n1373_o;
  wire n1375_o;
  wire n1376_o;
  wire n1378_o;
  wire n1379_o;
  wire n1381_o;
  wire n1382_o;
  wire n1384_o;
  wire n1386_o;
  wire n1388_o;
  wire n1389_o;
  wire n1391_o;
  wire n1393_o;
  wire n1394_o;
  wire n1396_o;
  wire n1397_o;
  wire n1399_o;
  wire n1400_o;
  wire n1402_o;
  wire n1403_o;
  wire n1405_o;
  wire n1406_o;
  wire n1408_o;
  wire n1409_o;
  wire n1411_o;
  wire n1412_o;
  wire n1414_o;
  wire n1415_o;
  wire n1417_o;
  wire n1418_o;
  wire n1420_o;
  wire n1421_o;
  wire n1423_o;
  wire n1425_o;
  wire n1427_o;
  wire n1428_o;
  wire n1430_o;
  wire n1431_o;
  wire n1433_o;
  wire n1434_o;
  wire n1436_o;
  wire n1437_o;
  wire n1439_o;
  wire n1440_o;
  wire n1442_o;
  wire n1443_o;
  wire n1445_o;
  wire n1446_o;
  wire n1448_o;
  wire n1450_o;
  wire n1451_o;
  wire n1453_o;
  wire n1455_o;
  wire n1456_o;
  wire n1458_o;
  wire n1460_o;
  wire n1461_o;
  wire n1463_o;
  wire n1464_o;
  wire n1466_o;
  wire n1467_o;
  wire n1469_o;
  wire n1470_o;
  wire n1472_o;
  wire n1473_o;
  wire n1475_o;
  wire n1476_o;
  wire n1478_o;
  wire n1479_o;
  wire n1481_o;
  wire n1483_o;
  wire n1485_o;
  wire n1487_o;
  wire n1488_o;
  wire n1490_o;
  wire n1491_o;
  wire n1493_o;
  wire n1494_o;
  wire n1496_o;
  wire n1498_o;
  wire n1500_o;
  wire n1501_o;
  wire n1503_o;
  wire n1505_o;
  wire n1507_o;
  wire n1509_o;
  wire n1510_o;
  wire n1512_o;
  wire n1513_o;
  wire n1515_o;
  wire n1516_o;
  wire n1518_o;
  wire n1519_o;
  wire n1521_o;
  wire n1522_o;
  wire n1524_o;
  wire n1525_o;
  wire n1527_o;
  wire n1528_o;
  wire n1530_o;
  wire n1531_o;
  wire n1533_o;
  wire n1534_o;
  wire n1536_o;
  wire n1538_o;
  wire n1540_o;
  wire n1541_o;
  wire n1543_o;
  wire n1544_o;
  wire n1546_o;
  wire n1547_o;
  wire n1549_o;
  wire n1550_o;
  wire n1552_o;
  wire n1553_o;
  wire n1555_o;
  wire n1556_o;
  wire n1558_o;
  wire n1559_o;
  wire n1561_o;
  wire n1562_o;
  wire n1564_o;
  wire n1565_o;
  wire n1567_o;
  wire n1569_o;
  wire n1570_o;
  wire n1572_o;
  wire n1573_o;
  wire n1575_o;
  wire n1576_o;
  wire n1578_o;
  wire n1579_o;
  wire n1581_o;
  wire n1582_o;
  wire n1584_o;
  wire n1585_o;
  wire n1587_o;
  wire n1588_o;
  wire n1590_o;
  wire n1591_o;
  wire n1593_o;
  wire n1594_o;
  wire n1596_o;
  wire n1598_o;
  wire n1599_o;
  wire n1601_o;
  wire n1603_o;
  wire n1604_o;
  wire n1606_o;
  wire n1607_o;
  wire n1609_o;
  wire n1610_o;
  wire n1612_o;
  wire n1614_o;
  wire n1615_o;
  wire n1617_o;
  wire n1619_o;
  wire n1620_o;
  wire n1622_o;
  wire n1623_o;
  wire n1625_o;
  wire n1626_o;
  wire n1628_o;
  wire n1630_o;
  wire n1632_o;
  wire n1633_o;
  wire n1635_o;
  wire n1636_o;
  wire n1638_o;
  wire n1639_o;
  wire n1641_o;
  wire n1642_o;
  wire n1644_o;
  wire n1645_o;
  wire n1647_o;
  wire n1648_o;
  wire n1650_o;
  wire n1651_o;
  wire n1653_o;
  wire n1654_o;
  wire n1656_o;
  wire n1657_o;
  wire n1659_o;
  wire n1661_o;
  wire n1663_o;
  wire n1664_o;
  wire n1666_o;
  wire n1667_o;
  wire n1669_o;
  wire n1671_o;
  wire n1672_o;
  wire n1674_o;
  wire n1675_o;
  wire n1677_o;
  wire n1678_o;
  wire n1680_o;
  wire n1681_o;
  wire n1683_o;
  wire n1684_o;
  wire n1686_o;
  wire n1687_o;
  wire n1689_o;
  wire n1690_o;
  wire n1692_o;
  wire n1693_o;
  wire n1695_o;
  wire n1696_o;
  wire n1698_o;
  wire n1699_o;
  wire n1701_o;
  wire n1702_o;
  wire n1704_o;
  wire n1706_o;
  wire n1707_o;
  wire n1709_o;
  wire n1710_o;
  wire n1712_o;
  wire n1714_o;
  wire n1715_o;
  wire n1717_o;
  wire n1719_o;
  wire n1720_o;
  wire n1722_o;
  wire n1724_o;
  wire n1725_o;
  wire n1727_o;
  wire n1729_o;
  wire n1730_o;
  wire n1732_o;
  wire n1734_o;
  wire n1735_o;
  wire n1737_o;
  wire n1739_o;
  wire n1741_o;
  wire n1742_o;
  wire n1744_o;
  wire n1746_o;
  wire n1748_o;
  wire n1749_o;
  wire n1751_o;
  wire n1752_o;
  wire n1754_o;
  wire n1755_o;
  wire n1757_o;
  wire n1758_o;
  wire n1760_o;
  wire n1761_o;
  wire n1763_o;
  wire n1764_o;
  wire n1766_o;
  wire n1767_o;
  wire n1769_o;
  wire n1770_o;
  wire n1772_o;
  wire n1773_o;
  wire n1775_o;
  wire n1776_o;
  wire n1778_o;
  wire n1779_o;
  wire n1781_o;
  wire n1783_o;
  wire n1784_o;
  wire n1786_o;
  wire n1787_o;
  wire n1789_o;
  wire n1790_o;
  wire n1792_o;
  wire n1793_o;
  wire n1795_o;
  wire n1796_o;
  wire n1798_o;
  wire n1799_o;
  wire n1801_o;
  wire n1802_o;
  wire n1804_o;
  wire n1805_o;
  wire n1807_o;
  wire n1808_o;
  wire n1810_o;
  wire [56:0] n1811_o;
  reg [5:0] n1870_o;
  reg n1900_o;
  wire [6:0] n1904_o;
  wire n1906_o;
  wire [5:0] n1908_o;
  wire [7:0] n1910_o;
  wire [5:0] n1911_o;
  wire [7:0] n1912_o;
  wire [5:0] n1913_o;
  wire n1923_o;
  wire [5:0] n1925_o;
  wire [5:0] n1926_o;
  wire int_b_n1927;
  wire int_b_n1929;
  wire int_b_n1930;
  wire int_b_n1931;
  wire int_b_tf_o;
  wire int_b_ext_int_o;
  wire int_b_tim_int_o;
  wire int_b_int_pending_o;
  wire int_b_int_in_progress_o;
  wire n1941_o;
  wire n1942_o;
  wire n1943_o;
  wire n1946_o;
  wire n1947_o;
  wire n1948_o;
  wire n1949_o;
  wire n1950_o;
  wire n1953_o;
  wire n1954_o;
  wire n1957_o;
  wire n1959_o;
  wire n1962_o;
  wire n1964_o;
  wire n1966_o;
  wire n1968_o;
  wire n1970_o;
  wire n1971_o;
  wire n1972_o;
  wire n1975_o;
  wire n1978_o;
  wire n1980_o;
  wire n1982_o;
  wire n1984_o;
  wire n1985_o;
  wire n1986_o;
  wire n1987_o;
  wire n1988_o;
  wire n1991_o;
  wire n1993_o;
  wire n1996_o;
  wire n1998_o;
  wire n1999_o;
  wire n2000_o;
  wire n2001_o;
  wire n2002_o;
  wire n2005_o;
  wire n2008_o;
  wire n2011_o;
  wire n2013_o;
  wire n2014_o;
  wire n2015_o;
  wire n2016_o;
  wire n2017_o;
  wire n2018_o;
  wire n2019_o;
  wire n2022_o;
  wire n2024_o;
  wire [4:0] n2025_o;
  reg n2027_o;
  reg n2030_o;
  reg n2033_o;
  reg n2036_o;
  reg n2039_o;
  reg n2042_o;
  reg n2045_o;
  reg n2048_o;
  reg n2051_o;
  wire n2058_o;
  wire n2059_o;
  wire n2061_o;
  wire n2062_o;
  wire n2063_o;
  wire [2:0] n2064_o;
  wire n2065_o;
  wire [2:0] n2067_o;
  wire [2:0] n2068_o;
  localparam [7:0] n2069_o = 8'b00000000;
  wire [4:0] n2070_o;
  wire n2073_o;
  wire [7:0] n2075_o;
  localparam [7:0] n2076_o = 8'bX;
  wire [7:0] n2077_o;
  wire n2081_o;
  wire n2083_o;
  wire n2084_o;
  wire n2086_o;
  wire n2093_o;
  wire n2096_o;
  wire [1:0] n2099_o;
  wire n2101_o;
  wire n2106_o;
  wire n2110_o;
  wire n2113_o;
  wire n2115_o;
  wire [2:0] n2116_o;
  reg n2119_o;
  reg n2122_o;
  reg n2125_o;
  reg n2126_o;
  reg n2129_o;
  reg [3:0] n2132_o;
  reg n2134_o;
  reg [1:0] n2136_o;
  reg n2138_o;
  reg n2141_o;
  reg n2144_o;
  wire n2146_o;
  wire n2148_o;
  wire n2152_o;
  wire n2155_o;
  wire n2157_o;
  wire [1:0] n2158_o;
  reg n2161_o;
  reg n2164_o;
  reg n2167_o;
  reg [3:0] n2170_o;
  reg n2172_o;
  reg n2174_o;
  reg n2177_o;
  reg n2180_o;
  wire n2182_o;
  wire n2184_o;
  wire n2186_o;
  wire [3:0] n2188_o;
  wire n2190_o;
  wire n2192_o;
  wire n2194_o;
  wire n2196_o;
  wire n2198_o;
  wire n2199_o;
  wire n2200_o;
  wire n2202_o;
  wire n2209_o;
  wire n2212_o;
  wire [1:0] n2215_o;
  wire n2217_o;
  wire n2222_o;
  wire n2227_o;
  wire [2:0] n2228_o;
  reg n2231_o;
  reg n2234_o;
  reg n2237_o;
  reg n2238_o;
  reg n2241_o;
  reg [3:0] n2244_o;
  reg [1:0] n2246_o;
  wire n2248_o;
  wire n2250_o;
  wire n2255_o;
  wire [1:0] n2256_o;
  reg n2259_o;
  reg n2262_o;
  reg n2265_o;
  reg [3:0] n2268_o;
  wire n2270_o;
  wire n2272_o;
  wire n2274_o;
  wire [3:0] n2276_o;
  wire n2278_o;
  wire n2279_o;
  wire n2281_o;
  wire [1:0] n2282_o;
  wire n2284_o;
  wire n2285_o;
  wire n2286_o;
  wire n2289_o;
  wire n2292_o;
  wire n2295_o;
  wire n2298_o;
  wire n2300_o;
  wire n2302_o;
  wire n2304_o;
  wire n2306_o;
  wire n2309_o;
  wire n2312_o;
  wire n2314_o;
  wire n2316_o;
  wire n2318_o;
  wire n2320_o;
  wire n2322_o;
  wire n2324_o;
  wire n2326_o;
  wire [1:0] n2327_o;
  wire n2329_o;
  wire n2330_o;
  wire n2331_o;
  wire n2334_o;
  wire n2337_o;
  wire n2340_o;
  wire n2342_o;
  wire n2344_o;
  wire n2346_o;
  wire [2:0] n2347_o;
  reg n2351_o;
  reg n2355_o;
  reg n2357_o;
  reg n2359_o;
  reg n2361_o;
  reg [3:0] n2364_o;
  wire n2366_o;
  wire n2368_o;
  wire n2370_o;
  wire n2372_o;
  wire n2374_o;
  wire n2376_o;
  wire n2378_o;
  wire n2380_o;
  wire [3:0] n2382_o;
  wire n2384_o;
  wire n2386_o;
  wire n2388_o;
  wire n2390_o;
  wire n2391_o;
  wire n2392_o;
  wire n2395_o;
  wire n2397_o;
  wire n2399_o;
  wire n2401_o;
  wire [2:0] n2402_o;
  reg n2405_o;
  reg n2408_o;
  reg n2411_o;
  reg n2414_o;
  reg n2417_o;
  reg [1:0] n2421_o;
  reg n2424_o;
  reg n2426_o;
  reg n2430_o;
  localparam [7:0] n2432_o = 8'b00000000;
  wire n2435_o;
  wire n2436_o;
  wire [4:0] n2437_o;
  wire [7:0] n2438_o;
  wire [7:0] n2439_o;
  wire n2441_o;
  wire n2443_o;
  wire n2444_o;
  wire [4:0] n2446_o;
  wire [2:0] n2447_o;
  wire [7:0] n2448_o;
  wire [7:0] n2450_o;
  wire n2453_o;
  wire n2455_o;
  wire [1:0] n2456_o;
  reg n2459_o;
  reg n2462_o;
  reg n2465_o;
  reg [7:0] n2466_o;
  reg n2468_o;
  reg n2470_o;
  wire n2471_o;
  wire n2473_o;
  wire n2475_o;
  wire n2477_o;
  wire n2479_o;
  wire n2481_o;
  wire n2483_o;
  wire [1:0] n2485_o;
  wire n2487_o;
  wire n2489_o;
  wire n2491_o;
  wire [7:0] n2492_o;
  wire n2493_o;
  wire n2495_o;
  wire n2497_o;
  wire n2499_o;
  wire n2501_o;
  wire n2504_o;
  wire n2507_o;
  wire [3:0] n2510_o;
  wire n2512_o;
  wire n2514_o;
  wire n2517_o;
  wire n2519_o;
  wire n2521_o;
  wire n2522_o;
  wire n2523_o;
  wire n2526_o;
  wire n2529_o;
  wire n2531_o;
  wire n2533_o;
  wire n2535_o;
  wire n2537_o;
  wire n2540_o;
  wire n2543_o;
  wire [3:0] n2546_o;
  wire n2548_o;
  wire n2550_o;
  wire n2551_o;
  wire n2553_o;
  wire n2556_o;
  wire n2558_o;
  wire n2560_o;
  wire n2561_o;
  wire n2562_o;
  wire n2563_o;
  wire n2565_o;
  wire n2568_o;
  wire n2571_o;
  wire n2573_o;
  wire n2575_o;
  wire n2577_o;
  wire n2579_o;
  wire n2581_o;
  wire n2582_o;
  wire n2585_o;
  wire n2588_o;
  wire n2590_o;
  wire [3:0] n2593_o;
  wire n2595_o;
  wire n2597_o;
  wire [2:0] n2598_o;
  reg n2601_o;
  reg n2603_o;
  reg n2606_o;
  reg [3:0] n2608_o;
  reg n2612_o;
  reg n2615_o;
  reg n2618_o;
  reg n2620_o;
  reg n2623_o;
  wire n2625_o;
  wire n2626_o;
  wire n2629_o;
  wire n2632_o;
  wire n2634_o;
  wire n2635_o;
  wire n2636_o;
  wire n2639_o;
  wire n2642_o;
  wire n2644_o;
  wire [1:0] n2645_o;
  reg n2647_o;
  reg n2649_o;
  reg n2652_o;
  reg n2654_o;
  reg [3:0] n2657_o;
  reg n2659_o;
  wire n2661_o;
  wire n2663_o;
  wire n2664_o;
  wire n2667_o;
  wire n2670_o;
  wire n2672_o;
  wire n2674_o;
  wire n2676_o;
  wire n2678_o;
  wire n2679_o;
  wire n2682_o;
  wire n2685_o;
  wire n2687_o;
  wire n2689_o;
  wire n2691_o;
  wire n2692_o;
  wire n2694_o;
  wire n2697_o;
  wire [1:0] n2698_o;
  reg n2701_o;
  reg n2704_o;
  reg n2707_o;
  reg [3:0] n2710_o;
  reg n2713_o;
  reg [3:0] n2716_o;
  wire n2717_o;
  reg n2718_o;
  reg n2721_o;
  wire n2723_o;
  wire n2724_o;
  wire n2730_o;
  wire n2733_o;
  wire n2735_o;
  wire n2737_o;
  wire n2739_o;
  wire n2741_o;
  wire [3:0] n2743_o;
  wire n2745_o;
  wire [3:0] n2747_o;
  wire n2748_o;
  wire n2749_o;
  wire n2751_o;
  wire n2753_o;
  wire n2755_o;
  wire n2757_o;
  wire n2760_o;
  wire n2762_o;
  wire n2764_o;
  wire n2765_o;
  wire n2766_o;
  wire n2767_o;
  wire n2770_o;
  wire n2773_o;
  wire n2776_o;
  wire n2778_o;
  wire n2780_o;
  wire n2782_o;
  wire n2784_o;
  wire n2785_o;
  wire n2788_o;
  wire n2791_o;
  wire n2793_o;
  wire n2794_o;
  wire n2795_o;
  wire n2797_o;
  wire n2804_o;
  wire n2807_o;
  wire [1:0] n2810_o;
  wire n2812_o;
  wire [1:0] n2813_o;
  wire n2815_o;
  wire n2818_o;
  wire n2821_o;
  wire n2823_o;
  wire [1:0] n2824_o;
  wire n2826_o;
  wire n2829_o;
  wire n2832_o;
  wire n2834_o;
  wire [2:0] n2835_o;
  reg n2837_o;
  reg n2839_o;
  reg n2842_o;
  reg n2843_o;
  reg n2845_o;
  reg [3:0] n2848_o;
  reg [1:0] n2850_o;
  reg n2852_o;
  wire n2854_o;
  wire n2855_o;
  wire n2857_o;
  wire n2860_o;
  wire n2863_o;
  wire n2865_o;
  wire n2866_o;
  wire n2872_o;
  wire n2875_o;
  wire n2877_o;
  wire n2879_o;
  wire n2881_o;
  wire n2883_o;
  wire n2885_o;
  wire n2886_o;
  wire n2888_o;
  wire n2889_o;
  wire n2892_o;
  wire n2893_o;
  wire n2894_o;
  wire n2896_o;
  wire n2897_o;
  wire n2903_o;
  wire n2906_o;
  wire n2908_o;
  wire n2910_o;
  wire n2912_o;
  wire n2914_o;
  wire n2916_o;
  wire n2917_o;
  wire n2919_o;
  wire n2920_o;
  wire [3:0] n2923_o;
  wire n2926_o;
  wire [3:0] n2928_o;
  wire n2930_o;
  wire n2931_o;
  wire n2937_o;
  wire n2940_o;
  wire n2942_o;
  wire n2944_o;
  wire [3:0] n2946_o;
  wire n2948_o;
  wire n2950_o;
  wire n2952_o;
  wire [4:0] n2954_o;
  wire [2:0] n2955_o;
  wire [7:0] n2956_o;
  wire n2958_o;
  wire [1:0] n2959_o;
  reg n2962_o;
  reg n2965_o;
  reg n2968_o;
  reg [7:0] n2969_o;
  reg n2971_o;
  wire n2973_o;
  wire n2975_o;
  wire n2977_o;
  wire [7:0] n2978_o;
  wire n2979_o;
  wire n2981_o;
  wire n2982_o;
  wire n2984_o;
  wire n2987_o;
  wire [1:0] n2990_o;
  wire n2992_o;
  wire n2995_o;
  wire n2998_o;
  wire n3000_o;
  wire n3002_o;
  wire [1:0] n3004_o;
  wire n3006_o;
  wire n3008_o;
  wire n3009_o;
  wire n3011_o;
  wire n3014_o;
  wire n3016_o;
  wire n3017_o;
  wire n3023_o;
  wire n3026_o;
  wire n3028_o;
  wire n3030_o;
  wire n3032_o;
  wire n3034_o;
  wire n3035_o;
  wire n3036_o;
  wire [3:0] n3039_o;
  wire n3040_o;
  wire n3042_o;
  wire n3043_o;
  wire n3046_o;
  wire n3047_o;
  wire n3048_o;
  wire n3050_o;
  wire n3051_o;
  wire n3057_o;
  wire n3060_o;
  wire n3062_o;
  wire n3064_o;
  wire n3066_o;
  wire n3068_o;
  wire n3070_o;
  wire n3071_o;
  wire n3073_o;
  wire n3076_o;
  wire n3079_o;
  wire n3081_o;
  wire n3082_o;
  wire n3088_o;
  wire n3091_o;
  wire n3093_o;
  wire n3095_o;
  wire n3097_o;
  wire n3099_o;
  wire n3101_o;
  wire n3102_o;
  wire n3104_o;
  wire n3105_o;
  wire n3108_o;
  wire n3111_o;
  wire n3112_o;
  wire n3113_o;
  wire n3115_o;
  wire n3116_o;
  wire n3122_o;
  wire n3125_o;
  wire n3127_o;
  wire n3129_o;
  wire n3131_o;
  wire n3133_o;
  wire n3135_o;
  wire n3137_o;
  wire n3139_o;
  wire n3140_o;
  wire n3143_o;
  wire n3145_o;
  wire n3146_o;
  wire n3147_o;
  wire n3149_o;
  wire n3156_o;
  wire n3159_o;
  wire [1:0] n3162_o;
  wire n3164_o;
  wire n3169_o;
  wire [1:0] n3170_o;
  reg n3173_o;
  reg n3176_o;
  reg n3177_o;
  reg n3180_o;
  reg [1:0] n3182_o;
  wire n3184_o;
  wire n3186_o;
  wire n3189_o;
  wire n3192_o;
  wire n3195_o;
  wire n3197_o;
  wire n3199_o;
  wire n3202_o;
  wire n3205_o;
  wire n3208_o;
  wire n3210_o;
  wire n3211_o;
  wire n3212_o;
  wire n3214_o;
  wire n3221_o;
  wire n3224_o;
  wire [1:0] n3227_o;
  wire n3229_o;
  wire n3231_o;
  wire [1:0] n3232_o;
  reg n3235_o;
  reg n3236_o;
  reg n3238_o;
  reg [1:0] n3240_o;
  reg n3243_o;
  wire n3245_o;
  wire n3246_o;
  wire n3248_o;
  wire n3249_o;
  wire n3250_o;
  wire n3251_o;
  wire n3253_o;
  wire n3260_o;
  wire n3263_o;
  wire [1:0] n3266_o;
  wire n3267_o;
  wire n3269_o;
  wire [1:0] n3271_o;
  wire n3273_o;
  wire n3274_o;
  wire n3277_o;
  wire n3279_o;
  wire n3281_o;
  wire n3282_o;
  wire n3285_o;
  wire n3288_o;
  wire n3291_o;
  wire n3294_o;
  wire n3296_o;
  wire n3298_o;
  wire n3300_o;
  wire n3302_o;
  wire n3304_o;
  wire n3305_o;
  wire [1:0] n3307_o;
  wire [3:0] n3308_o;
  wire n3311_o;
  wire n3314_o;
  wire n3317_o;
  wire [2:0] n3318_o;
  wire [1:0] n3319_o;
  wire [1:0] n3320_o;
  wire [1:0] n3321_o;
  reg [1:0] n3322_o;
  wire n3324_o;
  wire n3326_o;
  wire n3328_o;
  wire [2:0] n3329_o;
  reg n3332_o;
  reg n3336_o;
  wire [1:0] n3337_o;
  wire [1:0] n3338_o;
  wire [1:0] n3339_o;
  reg [1:0] n3340_o;
  wire [1:0] n3341_o;
  wire [1:0] n3342_o;
  wire [1:0] n3343_o;
  reg [1:0] n3344_o;
  wire [3:0] n3345_o;
  wire [3:0] n3346_o;
  wire [3:0] n3347_o;
  reg [3:0] n3348_o;
  reg n3350_o;
  reg n3354_o;
  wire n3356_o;
  wire n3358_o;
  wire n3359_o;
  wire n3362_o;
  wire n3364_o;
  wire n3366_o;
  wire [7:0] n3367_o;
  wire [7:0] n3368_o;
  wire n3369_o;
  wire n3370_o;
  wire n3372_o;
  wire n3373_o;
  wire [1:0] n3374_o;
  wire [7:0] n3376_o;
  wire n3378_o;
  wire n3381_o;
  wire n3383_o;
  wire [2:0] n3384_o;
  reg n3388_o;
  wire [3:0] n3389_o;
  wire [3:0] n3390_o;
  wire [3:0] n3391_o;
  wire [3:0] n3392_o;
  reg [3:0] n3393_o;
  wire [3:0] n3394_o;
  wire [3:0] n3395_o;
  wire [3:0] n3396_o;
  wire [3:0] n3397_o;
  reg [3:0] n3398_o;
  reg n3401_o;
  reg n3405_o;
  wire n3407_o;
  wire n3409_o;
  wire [1:0] n3410_o;
  reg n3413_o;
  reg n3416_o;
  reg n3419_o;
  reg n3423_o;
  wire n3425_o;
  wire n3427_o;
  wire n3429_o;
  wire n3431_o;
  wire [7:0] n3432_o;
  wire [7:0] n3433_o;
  wire n3434_o;
  wire n3435_o;
  wire n3437_o;
  wire n3438_o;
  wire n3440_o;
  wire n3441_o;
  wire n3442_o;
  wire [1:0] n3445_o;
  wire n3448_o;
  wire [1:0] n3450_o;
  wire n3452_o;
  wire n3455_o;
  wire n3458_o;
  wire n3460_o;
  wire n3462_o;
  wire [1:0] n3464_o;
  wire n3466_o;
  wire n3468_o;
  wire n3469_o;
  wire n3470_o;
  wire n3473_o;
  wire n3476_o;
  wire n3477_o;
  wire n3479_o;
  wire n3480_o;
  wire n3483_o;
  wire n3486_o;
  wire n3488_o;
  wire [1:0] n3489_o;
  reg n3491_o;
  reg n3494_o;
  reg n3497_o;
  wire n3499_o;
  wire n3500_o;
  wire n3501_o;
  wire n3504_o;
  wire n3507_o;
  wire n3510_o;
  wire n3513_o;
  wire n3515_o;
  wire n3517_o;
  wire n3519_o;
  wire n3521_o;
  wire n3523_o;
  wire n3524_o;
  wire n3525_o;
  wire n3527_o;
  wire n3529_o;
  wire n3532_o;
  wire n3534_o;
  wire n3536_o;
  wire n3537_o;
  wire n3538_o;
  wire n3540_o;
  wire n3547_o;
  wire n3550_o;
  wire [1:0] n3553_o;
  wire n3555_o;
  wire n3560_o;
  wire n3565_o;
  wire [2:0] n3566_o;
  reg n3569_o;
  reg n3572_o;
  reg n3575_o;
  reg n3576_o;
  reg n3579_o;
  reg [3:0] n3582_o;
  reg [1:0] n3584_o;
  wire n3586_o;
  wire n3588_o;
  wire n3593_o;
  wire [1:0] n3594_o;
  reg n3597_o;
  reg n3600_o;
  reg n3603_o;
  reg [3:0] n3606_o;
  wire n3608_o;
  wire n3610_o;
  wire n3612_o;
  wire [3:0] n3614_o;
  wire n3616_o;
  wire n3617_o;
  wire n3619_o;
  wire [1:0] n3620_o;
  wire n3622_o;
  wire n3623_o;
  wire n3624_o;
  wire n3627_o;
  wire n3630_o;
  wire n3633_o;
  wire n3636_o;
  wire n3638_o;
  wire n3640_o;
  wire n3642_o;
  wire n3644_o;
  wire n3647_o;
  wire n3650_o;
  wire n3652_o;
  wire n3654_o;
  wire n3656_o;
  wire n3658_o;
  wire n3660_o;
  wire n3662_o;
  wire n3664_o;
  wire [1:0] n3665_o;
  wire n3667_o;
  wire n3668_o;
  wire n3669_o;
  wire n3672_o;
  wire n3675_o;
  wire n3678_o;
  wire n3680_o;
  wire n3682_o;
  wire n3684_o;
  wire [2:0] n3685_o;
  reg n3689_o;
  reg n3693_o;
  reg n3695_o;
  reg n3697_o;
  reg n3699_o;
  reg [3:0] n3702_o;
  wire n3704_o;
  wire n3706_o;
  wire n3708_o;
  wire n3710_o;
  wire n3712_o;
  wire n3714_o;
  wire n3716_o;
  wire n3718_o;
  wire [3:0] n3720_o;
  wire n3722_o;
  wire n3724_o;
  wire n3726_o;
  wire n3728_o;
  wire n3729_o;
  wire n3730_o;
  wire n3733_o;
  wire n3734_o;
  wire n3736_o;
  wire n3737_o;
  wire n3738_o;
  wire n3739_o;
  wire n3740_o;
  wire n3743_o;
  wire n3746_o;
  wire n3749_o;
  wire n3751_o;
  wire n3753_o;
  wire n3756_o;
  wire n3758_o;
  wire n3760_o;
  wire n3762_o;
  wire n3764_o;
  wire n3765_o;
  wire n3767_o;
  wire n3769_o;
  wire n3771_o;
  wire [2:0] n3772_o;
  reg n3775_o;
  reg n3778_o;
  reg n3781_o;
  reg n3784_o;
  reg [1:0] n3788_o;
  reg n3791_o;
  wire n3792_o;
  wire n3795_o;
  wire n3798_o;
  wire n3800_o;
  wire n3802_o;
  wire [1:0] n3803_o;
  reg n3806_o;
  reg n3809_o;
  reg n3811_o;
  reg n3814_o;
  reg n3816_o;
  wire n3817_o;
  wire n3818_o;
  wire n3820_o;
  wire n3822_o;
  wire n3824_o;
  wire n3826_o;
  wire [1:0] n3828_o;
  wire n3830_o;
  wire n3832_o;
  wire n3834_o;
  wire n3836_o;
  wire n3838_o;
  wire n3839_o;
  wire n3842_o;
  wire n3844_o;
  wire n3847_o;
  wire n3850_o;
  wire n3853_o;
  wire [3:0] n3856_o;
  wire n3858_o;
  wire n3860_o;
  wire n3862_o;
  wire n3864_o;
  wire n3866_o;
  wire n3867_o;
  wire n3868_o;
  wire n3871_o;
  wire n3873_o;
  wire n3876_o;
  wire n3879_o;
  wire n3882_o;
  wire [3:0] n3885_o;
  wire n3887_o;
  wire n3889_o;
  wire n3891_o;
  wire n3893_o;
  wire n3895_o;
  wire n3896_o;
  wire n3899_o;
  wire n3902_o;
  wire n3904_o;
  wire n3906_o;
  wire n3908_o;
  wire n3910_o;
  wire n3911_o;
  wire n3913_o;
  wire n3916_o;
  wire n3918_o;
  wire n3920_o;
  wire n3923_o;
  wire n3925_o;
  wire n3927_o;
  wire n3928_o;
  wire n3931_o;
  wire n3934_o;
  wire n3936_o;
  wire n3938_o;
  wire n3940_o;
  wire n3942_o;
  wire n3945_o;
  wire n3948_o;
  wire n3950_o;
  wire n3951_o;
  wire n3952_o;
  wire n3954_o;
  wire n3961_o;
  wire n3964_o;
  wire [1:0] n3967_o;
  wire n3969_o;
  wire n3970_o;
  wire n3973_o;
  wire n3975_o;
  wire n3976_o;
  wire [3:0] n3979_o;
  wire n3981_o;
  wire [2:0] n3982_o;
  reg n3985_o;
  reg n3988_o;
  reg n3991_o;
  reg n3992_o;
  reg n3995_o;
  reg [3:0] n3997_o;
  reg n3999_o;
  reg [1:0] n4001_o;
  reg n4004_o;
  wire n4006_o;
  wire n4007_o;
  wire n4008_o;
  wire n4010_o;
  wire n4017_o;
  wire n4020_o;
  wire [1:0] n4023_o;
  wire n4025_o;
  wire n4030_o;
  wire n4035_o;
  wire [2:0] n4036_o;
  reg n4039_o;
  reg n4042_o;
  reg n4045_o;
  reg n4046_o;
  reg n4049_o;
  reg [3:0] n4052_o;
  reg [1:0] n4054_o;
  wire n4056_o;
  wire n4058_o;
  wire n4063_o;
  wire [1:0] n4064_o;
  reg n4067_o;
  reg n4070_o;
  reg n4073_o;
  reg [3:0] n4076_o;
  wire n4078_o;
  wire n4080_o;
  wire n4082_o;
  wire [3:0] n4084_o;
  wire n4086_o;
  wire [56:0] n4087_o;
  reg n4089_o;
  reg n4092_o;
  reg n4095_o;
  reg n4098_o;
  reg n4101_o;
  reg n4103_o;
  reg n4105_o;
  reg n4108_o;
  reg n4111_o;
  reg n4114_o;
  reg n4117_o;
  reg n4120_o;
  reg n4123_o;
  reg n4126_o;
  reg n4129_o;
  reg n4132_o;
  reg n4135_o;
  reg n4138_o;
  reg n4141_o;
  reg n4144_o;
  reg n4147_o;
  reg [3:0] n4151_o;
  reg n4154_o;
  reg n4157_o;
  reg n4160_o;
  reg n4163_o;
  reg n4166_o;
  reg n4170_o;
  reg n4175_o;
  reg n4179_o;
  reg n4182_o;
  reg n4185_o;
  reg [3:0] n4193_o;
  wire n4195_o;
  reg n4196_o;
  wire [1:0] n4197_o;
  reg [1:0] n4199_o;
  reg n4202_o;
  reg n4205_o;
  reg [1:0] n4208_o;
  reg n4211_o;
  reg n4214_o;
  reg n4217_o;
  reg n4220_o;
  reg n4223_o;
  reg n4226_o;
  reg n4229_o;
  reg n4232_o;
  reg n4235_o;
  reg n4238_o;
  reg n4241_o;
  reg n4244_o;
  reg n4267_o;
  reg n4270_o;
  reg n4273_o;
  reg n4276_o;
  reg n4279_o;
  reg n4282_o;
  reg n4285_o;
  reg n4288_o;
  reg n4291_o;
  reg [7:0] n4293_o;
  reg n4294_o;
  reg n4296_o;
  reg n4299_o;
  reg n4302_o;
  reg n4305_o;
  reg n4308_o;
  reg n4311_o;
  reg n4314_o;
  reg n4317_o;
  reg n4320_o;
  reg n4323_o;
  reg n4326_o;
  wire n4330_o;
  wire n4333_o;
  wire n4335_o;
  wire n4337_o;
  wire n4338_o;
  wire n4339_o;
  wire n4341_o;
  wire n4343_o;
  wire n4345_o;
  wire n4351_o;
  wire [7:0] n4365_o;
  wire n4367_o;
  wire n4368_o;
  wire n4369_o;
  wire n4370_o;
  wire [7:0] n4371_o;
  reg [7:0] n4372_q;
  wire n4373_o;
  reg n4374_q;
  wire n4375_o;
  reg n4376_q;
  wire n4377_o;
  reg n4378_q;
  wire n4379_o;
  reg n4380_q;
  wire [5:0] n4381_o;
  reg [5:0] n4382_q;
  wire [2:0] n4383_o;
  assign t0_dir_o = t0_dir_q;
  assign data_o = n4365_o;
  assign alu_write_accu_o = n4089_o;
  assign alu_write_shadow_o = n4092_o;
  assign alu_write_temp_reg_o = n4095_o;
  assign alu_read_alu_o = n4098_o;
  assign bus_write_bus_o = n4101_o;
  assign bus_read_bus_o = n4370_o;
  assign dm_write_dmem_addr_o = n4103_o;
  assign dm_write_dmem_o = n4367_o;
  assign dm_read_dmem_o = n4105_o;
  assign p1_write_p1_o = n4108_o;
  assign p1_read_p1_o = n4111_o;
  assign p2_write_p2_o = n4114_o;
  assign p2_write_exp_o = n4117_o;
  assign p2_read_p2_o = n4120_o;
  assign p2_read_exp_o = n4123_o;
  assign pm_write_pcl_o = n4126_o;
  assign pm_read_pcl_o = n4129_o;
  assign pm_write_pch_o = n4132_o;
  assign pm_read_pch_o = n4135_o;
  assign pm_read_pmem_o = n2027_o;
  assign psw_read_psw_o = n4138_o;
  assign psw_read_sp_o = n4141_o;
  assign psw_write_psw_o = n4144_o;
  assign psw_write_sp_o = n4147_o;
  assign alu_op_o = n4151_o;
  assign alu_use_carry_o = n4154_o;
  assign alu_da_high_o = n4157_o;
  assign alu_accu_low_o = n4160_o;
  assign alu_p06_temp_reg_o = n4163_o;
  assign alu_p60_temp_reg_o = n4166_o;
  assign bus_output_pcl_o = n2030_o;
  assign bus_bidir_bus_o = n4170_o;
  assign clk_multi_cycle_o = opc_multi_cycle_s;
  assign clk_assert_psen_o = n2033_o;
  assign clk_assert_prog_o = n4175_o;
  assign clk_assert_rd_o = n4179_o;
  assign clk_assert_wr_o = n4182_o;
  assign cnd_compute_take_o = n4185_o;
  assign cnd_branch_cond_o = n4193_o;
  assign cnd_comp_value_o = n4383_o;
  assign cnd_f1_o = f1_q;
  assign cnd_tf_o = tf_s;
  assign dm_addr_type_o = n4199_o;
  assign p1_read_reg_o = n4202_o;
  assign p2_read_reg_o = n4205_o;
  assign p2_output_pch_o = n2036_o;
  assign pm_inc_pc_o = n4368_o;
  assign pm_write_pmem_addr_o = n4369_o;
  assign pm_addr_type_o = n4208_o;
  assign psw_special_data_o = n4211_o;
  assign psw_inc_stackp_o = n4214_o;
  assign psw_dec_stackp_o = n4217_o;
  assign psw_write_carry_o = n4220_o;
  assign psw_write_aux_carry_o = n4223_o;
  assign psw_write_f0_o = n4226_o;
  assign psw_write_bs_o = n4229_o;
  assign tim_read_timer_o = n4232_o;
  assign tim_write_timer_o = n4235_o;
  assign tim_start_t_o = n4238_o;
  assign tim_start_cnt_o = n4241_o;
  assign tim_stop_tcnt_o = n4244_o;
  /* decoder.vhd:179:10  */
  assign opc_multi_cycle_s = n1923_o; // (signal)
  /* decoder.vhd:180:10  */
  assign opc_read_bus_s = n2039_o; // (signal)
  /* decoder.vhd:181:10  */
  assign opc_inj_int_s = n2042_o; // (signal)
  /* decoder.vhd:182:10  */
  assign opc_opcode_q = n4372_q; // (signal)
  /* decoder.vhd:183:10  */
  assign opc_mnemonic_s = n1925_o; // (signal)
  /* decoder.vhd:184:10  */
  assign last_cycle_s = n1943_o; // (signal)
  /* decoder.vhd:187:10  */
  assign assert_psen_s = n4267_o; // (signal)
  /* decoder.vhd:190:10  */
  assign branch_taken_s = n4270_o; // (signal)

  always @(posedge clk_i)
  begin
    //if(en_clk_i && ale_i && cnd_take_branch_i) $display("cnd_take_branch_i branch_taken_s=%b opc_opcode_q=%x", branch_taken_s, opc_opcode_q);
  end


  /* decoder.vhd:191:10  */
  assign branch_taken_q = n4374_q; // (signal)
  /* decoder.vhd:192:10  */
  assign pm_inc_pc_s = n2045_o; // (signal)
  /* decoder.vhd:193:10  */
  assign pm_write_pmem_addr_s = n2048_o; // (signal)
  /* decoder.vhd:195:10  */
  assign add_inc_pc_s = n4273_o; // (signal)
  /* decoder.vhd:197:10  */
  assign add_write_pmem_addr_s = n4276_o; // (signal)
  /* decoder.vhd:200:10  */
  assign clear_f1_s = n4279_o; // (signal)
  /* decoder.vhd:201:10  */
  assign cpl_f1_s = n4282_o; // (signal)
  /* decoder.vhd:202:10  */
  assign f1_q = n4376_q; // (signal)
  /* decoder.vhd:204:10  */
  assign clear_mb_s = n4285_o; // (signal)
  /* decoder.vhd:205:10  */
  assign set_mb_s = n4288_o; // (signal)
  /* decoder.vhd:206:10  */
  assign mb_q = n4378_q; // (signal)
  /* decoder.vhd:209:10  */
  assign ent0_clk_s = n4291_o; // (signal)
  /* decoder.vhd:210:10  */
  assign t0_dir_q = n4380_q; // (signal)
  /* decoder.vhd:212:10  */
  assign data_s = n4293_o; // (signal)
  /* decoder.vhd:213:10  */
  assign read_dec_s = n4294_o; // (signal)
  /* decoder.vhd:215:10  */
  assign tf_s = int_b_n1927; // (signal)
  /* decoder.vhd:217:10  */
  assign bus_read_bus_s = n2051_o; // (signal)
  /* decoder.vhd:218:10  */
  assign add_read_bus_s = n4296_o; // (signal)
  /* decoder.vhd:220:10  */
  assign dm_write_dmem_s = n4299_o; // (signal)
  /* decoder.vhd:222:10  */
  assign p2_output_exp_s = n4302_o; // (signal)
  /* decoder.vhd:224:10  */
  assign movx_first_cycle_s = n4305_o; // (signal)
  /* decoder.vhd:227:10  */
  assign jtf_executed_s = n4308_o; // (signal)
  /* decoder.vhd:228:10  */
  assign en_tcnti_s = n4311_o; // (signal)
  /* decoder.vhd:229:10  */
  assign dis_tcnti_s = n4314_o; // (signal)
  /* decoder.vhd:230:10  */
  assign en_i_s = n4317_o; // (signal)
  /* decoder.vhd:231:10  */
  assign dis_i_s = n4320_o; // (signal)
  /* decoder.vhd:232:10  */
  assign tim_int_s = int_b_n1929; // (signal)
  /* decoder.vhd:233:10  */
  assign retr_executed_s = n4323_o; // (signal)
  /* decoder.vhd:234:10  */
  assign int_executed_s = n4326_o; // (signal)
  /* decoder.vhd:235:10  */
  assign int_pending_s = int_b_n1930; // (signal)
  /* decoder.vhd:236:10  */
  assign int_in_progress_s = int_b_n1931; // (signal)
  /* decoder.vhd:239:10  */
  assign mnemonic_rec_s = n1904_o; // (signal)
  /* decoder.vhd:240:10  */
  assign mnemonic_q = n4382_q; // (signal)
  /* decoder_pack-p.vhd:105:7  */
  assign n1179_o = opc_opcode_q == 8'b01101000;
  /* decoder_pack-p.vhd:105:23  */
  assign n1181_o = opc_opcode_q == 8'b01101001;
  /* decoder_pack-p.vhd:105:23  */
  assign n1182_o = n1179_o | n1181_o;
  /* decoder_pack-p.vhd:105:36  */
  assign n1184_o = opc_opcode_q == 8'b01101010;
  /* decoder_pack-p.vhd:105:36  */
  assign n1185_o = n1182_o | n1184_o;
  /* decoder_pack-p.vhd:105:49  */
  assign n1187_o = opc_opcode_q == 8'b01101011;
  /* decoder_pack-p.vhd:105:49  */
  assign n1188_o = n1185_o | n1187_o;
  /* decoder_pack-p.vhd:105:62  */
  assign n1190_o = opc_opcode_q == 8'b01101100;
  /* decoder_pack-p.vhd:105:62  */
  assign n1191_o = n1188_o | n1190_o;
  /* decoder_pack-p.vhd:106:23  */
  assign n1193_o = opc_opcode_q == 8'b01101101;
  /* decoder_pack-p.vhd:106:23  */
  assign n1194_o = n1191_o | n1193_o;
  /* decoder_pack-p.vhd:106:36  */
  assign n1196_o = opc_opcode_q == 8'b01101110;
  /* decoder_pack-p.vhd:106:36  */
  assign n1197_o = n1194_o | n1196_o;
  /* decoder_pack-p.vhd:106:49  */
  assign n1199_o = opc_opcode_q == 8'b01101111;
  /* decoder_pack-p.vhd:106:49  */
  assign n1200_o = n1197_o | n1199_o;
  /* decoder_pack-p.vhd:106:62  */
  assign n1202_o = opc_opcode_q == 8'b01100000;
  /* decoder_pack-p.vhd:106:62  */
  assign n1203_o = n1200_o | n1202_o;
  /* decoder_pack-p.vhd:107:23  */
  assign n1205_o = opc_opcode_q == 8'b01100001;
  /* decoder_pack-p.vhd:107:23  */
  assign n1206_o = n1203_o | n1205_o;
  /* decoder_pack-p.vhd:107:36  */
  assign n1208_o = opc_opcode_q == 8'b01111000;
  /* decoder_pack-p.vhd:107:36  */
  assign n1209_o = n1206_o | n1208_o;
  /* decoder_pack-p.vhd:108:23  */
  assign n1211_o = opc_opcode_q == 8'b01111001;
  /* decoder_pack-p.vhd:108:23  */
  assign n1212_o = n1209_o | n1211_o;
  /* decoder_pack-p.vhd:108:36  */
  assign n1214_o = opc_opcode_q == 8'b01111010;
  /* decoder_pack-p.vhd:108:36  */
  assign n1215_o = n1212_o | n1214_o;
  /* decoder_pack-p.vhd:108:49  */
  assign n1217_o = opc_opcode_q == 8'b01111011;
  /* decoder_pack-p.vhd:108:49  */
  assign n1218_o = n1215_o | n1217_o;
  /* decoder_pack-p.vhd:108:62  */
  assign n1220_o = opc_opcode_q == 8'b01111100;
  /* decoder_pack-p.vhd:108:62  */
  assign n1221_o = n1218_o | n1220_o;
  /* decoder_pack-p.vhd:109:23  */
  assign n1223_o = opc_opcode_q == 8'b01111101;
  /* decoder_pack-p.vhd:109:23  */
  assign n1224_o = n1221_o | n1223_o;
  /* decoder_pack-p.vhd:109:36  */
  assign n1226_o = opc_opcode_q == 8'b01111110;
  /* decoder_pack-p.vhd:109:36  */
  assign n1227_o = n1224_o | n1226_o;
  /* decoder_pack-p.vhd:109:49  */
  assign n1229_o = opc_opcode_q == 8'b01111111;
  /* decoder_pack-p.vhd:109:49  */
  assign n1230_o = n1227_o | n1229_o;
  /* decoder_pack-p.vhd:109:62  */
  assign n1232_o = opc_opcode_q == 8'b01110000;
  /* decoder_pack-p.vhd:109:62  */
  assign n1233_o = n1230_o | n1232_o;
  /* decoder_pack-p.vhd:110:23  */
  assign n1235_o = opc_opcode_q == 8'b01110001;
  /* decoder_pack-p.vhd:110:23  */
  assign n1236_o = n1233_o | n1235_o;
  /* decoder_pack-p.vhd:114:7  */
  assign n1238_o = opc_opcode_q == 8'b00000011;
  /* decoder_pack-p.vhd:114:23  */
  assign n1240_o = opc_opcode_q == 8'b00010011;
  /* decoder_pack-p.vhd:114:23  */
  assign n1241_o = n1238_o | n1240_o;
  /* decoder_pack-p.vhd:120:7  */
  assign n1243_o = opc_opcode_q == 8'b01011000;
  /* decoder_pack-p.vhd:120:23  */
  assign n1245_o = opc_opcode_q == 8'b01011001;
  /* decoder_pack-p.vhd:120:23  */
  assign n1246_o = n1243_o | n1245_o;
  /* decoder_pack-p.vhd:120:36  */
  assign n1248_o = opc_opcode_q == 8'b01011010;
  /* decoder_pack-p.vhd:120:36  */
  assign n1249_o = n1246_o | n1248_o;
  /* decoder_pack-p.vhd:120:49  */
  assign n1251_o = opc_opcode_q == 8'b01011011;
  /* decoder_pack-p.vhd:120:49  */
  assign n1252_o = n1249_o | n1251_o;
  /* decoder_pack-p.vhd:120:62  */
  assign n1254_o = opc_opcode_q == 8'b01011100;
  /* decoder_pack-p.vhd:120:62  */
  assign n1255_o = n1252_o | n1254_o;
  /* decoder_pack-p.vhd:121:23  */
  assign n1257_o = opc_opcode_q == 8'b01011101;
  /* decoder_pack-p.vhd:121:23  */
  assign n1258_o = n1255_o | n1257_o;
  /* decoder_pack-p.vhd:121:36  */
  assign n1260_o = opc_opcode_q == 8'b01011110;
  /* decoder_pack-p.vhd:121:36  */
  assign n1261_o = n1258_o | n1260_o;
  /* decoder_pack-p.vhd:121:49  */
  assign n1263_o = opc_opcode_q == 8'b01011111;
  /* decoder_pack-p.vhd:121:49  */
  assign n1264_o = n1261_o | n1263_o;
  /* decoder_pack-p.vhd:121:62  */
  assign n1266_o = opc_opcode_q == 8'b01010000;
  /* decoder_pack-p.vhd:121:62  */
  assign n1267_o = n1264_o | n1266_o;
  /* decoder_pack-p.vhd:122:23  */
  assign n1269_o = opc_opcode_q == 8'b01010001;
  /* decoder_pack-p.vhd:122:23  */
  assign n1270_o = n1267_o | n1269_o;
  /* decoder_pack-p.vhd:126:7  */
  assign n1272_o = opc_opcode_q == 8'b01010011;
  /* decoder_pack-p.vhd:131:7  */
  assign n1274_o = opc_opcode_q == 8'b10011000;
  /* decoder_pack-p.vhd:131:23  */
  assign n1276_o = opc_opcode_q == 8'b10011001;
  /* decoder_pack-p.vhd:131:23  */
  assign n1277_o = n1274_o | n1276_o;
  /* decoder_pack-p.vhd:132:23  */
  assign n1279_o = opc_opcode_q == 8'b10011010;
  /* decoder_pack-p.vhd:132:23  */
  assign n1280_o = n1277_o | n1279_o;
  /* decoder_pack-p.vhd:137:7  */
  assign n1282_o = opc_opcode_q == 8'b00010100;
  /* decoder_pack-p.vhd:137:23  */
  assign n1284_o = opc_opcode_q == 8'b00110100;
  /* decoder_pack-p.vhd:137:23  */
  assign n1285_o = n1282_o | n1284_o;
  /* decoder_pack-p.vhd:137:36  */
  assign n1287_o = opc_opcode_q == 8'b01010100;
  /* decoder_pack-p.vhd:137:36  */
  assign n1288_o = n1285_o | n1287_o;
  /* decoder_pack-p.vhd:137:49  */
  assign n1290_o = opc_opcode_q == 8'b01110100;
  /* decoder_pack-p.vhd:137:49  */
  assign n1291_o = n1288_o | n1290_o;
  /* decoder_pack-p.vhd:137:62  */
  assign n1293_o = opc_opcode_q == 8'b10010100;
  /* decoder_pack-p.vhd:137:62  */
  assign n1294_o = n1291_o | n1293_o;
  /* decoder_pack-p.vhd:138:23  */
  assign n1296_o = opc_opcode_q == 8'b10110100;
  /* decoder_pack-p.vhd:138:23  */
  assign n1297_o = n1294_o | n1296_o;
  /* decoder_pack-p.vhd:138:36  */
  assign n1299_o = opc_opcode_q == 8'b11010100;
  /* decoder_pack-p.vhd:138:36  */
  assign n1300_o = n1297_o | n1299_o;
  /* decoder_pack-p.vhd:138:49  */
  assign n1302_o = opc_opcode_q == 8'b11110100;
  /* decoder_pack-p.vhd:138:49  */
  assign n1303_o = n1300_o | n1302_o;
  /* decoder_pack-p.vhd:143:7  */
  assign n1305_o = opc_opcode_q == 8'b00100111;
  /* decoder_pack-p.vhd:147:7  */
  assign n1307_o = opc_opcode_q == 8'b10010111;
  /* decoder_pack-p.vhd:151:7  */
  assign n1309_o = opc_opcode_q == 8'b10000101;
  /* decoder_pack-p.vhd:151:23  */
  assign n1311_o = opc_opcode_q == 8'b10100101;
  /* decoder_pack-p.vhd:151:23  */
  assign n1312_o = n1309_o | n1311_o;
  /* decoder_pack-p.vhd:156:7  */
  assign n1314_o = opc_opcode_q == 8'b00110111;
  /* decoder_pack-p.vhd:160:7  */
  assign n1316_o = opc_opcode_q == 8'b10100111;
  /* decoder_pack-p.vhd:164:7  */
  assign n1318_o = opc_opcode_q == 8'b10010101;
  /* decoder_pack-p.vhd:164:23  */
  assign n1320_o = opc_opcode_q == 8'b10110101;
  /* decoder_pack-p.vhd:164:23  */
  assign n1321_o = n1318_o | n1320_o;
  /* decoder_pack-p.vhd:169:7  */
  assign n1323_o = opc_opcode_q == 8'b01010111;
  /* decoder_pack-p.vhd:173:7  */
  assign n1325_o = opc_opcode_q == 8'b11001000;
  /* decoder_pack-p.vhd:173:23  */
  assign n1327_o = opc_opcode_q == 8'b11001001;
  /* decoder_pack-p.vhd:173:23  */
  assign n1328_o = n1325_o | n1327_o;
  /* decoder_pack-p.vhd:173:36  */
  assign n1330_o = opc_opcode_q == 8'b11001010;
  /* decoder_pack-p.vhd:173:36  */
  assign n1331_o = n1328_o | n1330_o;
  /* decoder_pack-p.vhd:173:49  */
  assign n1333_o = opc_opcode_q == 8'b11001011;
  /* decoder_pack-p.vhd:173:49  */
  assign n1334_o = n1331_o | n1333_o;
  /* decoder_pack-p.vhd:173:62  */
  assign n1336_o = opc_opcode_q == 8'b11001100;
  /* decoder_pack-p.vhd:173:62  */
  assign n1337_o = n1334_o | n1336_o;
  /* decoder_pack-p.vhd:174:23  */
  assign n1339_o = opc_opcode_q == 8'b11001101;
  /* decoder_pack-p.vhd:174:23  */
  assign n1340_o = n1337_o | n1339_o;
  /* decoder_pack-p.vhd:174:36  */
  assign n1342_o = opc_opcode_q == 8'b11001110;
  /* decoder_pack-p.vhd:174:36  */
  assign n1343_o = n1340_o | n1342_o;
  /* decoder_pack-p.vhd:174:49  */
  assign n1345_o = opc_opcode_q == 8'b11001111;
  /* decoder_pack-p.vhd:174:49  */
  assign n1346_o = n1343_o | n1345_o;
  /* decoder_pack-p.vhd:174:62  */
  assign n1348_o = opc_opcode_q == 8'b00000111;
  /* decoder_pack-p.vhd:174:62  */
  assign n1349_o = n1346_o | n1348_o;
  /* decoder_pack-p.vhd:179:7  */
  assign n1351_o = opc_opcode_q == 8'b00010101;
  /* decoder_pack-p.vhd:179:23  */
  assign n1353_o = opc_opcode_q == 8'b00000101;
  /* decoder_pack-p.vhd:179:23  */
  assign n1354_o = n1351_o | n1353_o;
  /* decoder_pack-p.vhd:184:7  */
  assign n1356_o = opc_opcode_q == 8'b00110101;
  /* decoder_pack-p.vhd:184:23  */
  assign n1358_o = opc_opcode_q == 8'b00100101;
  /* decoder_pack-p.vhd:184:23  */
  assign n1359_o = n1356_o | n1358_o;
  /* decoder_pack-p.vhd:189:7  */
  assign n1361_o = opc_opcode_q == 8'b11101000;
  /* decoder_pack-p.vhd:189:23  */
  assign n1363_o = opc_opcode_q == 8'b11101001;
  /* decoder_pack-p.vhd:189:23  */
  assign n1364_o = n1361_o | n1363_o;
  /* decoder_pack-p.vhd:189:36  */
  assign n1366_o = opc_opcode_q == 8'b11101010;
  /* decoder_pack-p.vhd:189:36  */
  assign n1367_o = n1364_o | n1366_o;
  /* decoder_pack-p.vhd:189:49  */
  assign n1369_o = opc_opcode_q == 8'b11101011;
  /* decoder_pack-p.vhd:189:49  */
  assign n1370_o = n1367_o | n1369_o;
  /* decoder_pack-p.vhd:189:62  */
  assign n1372_o = opc_opcode_q == 8'b11101100;
  /* decoder_pack-p.vhd:189:62  */
  assign n1373_o = n1370_o | n1372_o;
  /* decoder_pack-p.vhd:190:23  */
  assign n1375_o = opc_opcode_q == 8'b11101101;
  /* decoder_pack-p.vhd:190:23  */
  assign n1376_o = n1373_o | n1375_o;
  /* decoder_pack-p.vhd:190:36  */
  assign n1378_o = opc_opcode_q == 8'b11101110;
  /* decoder_pack-p.vhd:190:36  */
  assign n1379_o = n1376_o | n1378_o;
  /* decoder_pack-p.vhd:190:49  */
  assign n1381_o = opc_opcode_q == 8'b11101111;
  /* decoder_pack-p.vhd:190:49  */
  assign n1382_o = n1379_o | n1381_o;
  /* decoder_pack-p.vhd:195:7  */
  assign n1384_o = opc_opcode_q == 8'b01110101;
  /* decoder_pack-p.vhd:199:7  */
  assign n1386_o = opc_opcode_q == 8'b00001001;
  /* decoder_pack-p.vhd:199:23  */
  assign n1388_o = opc_opcode_q == 8'b00001010;
  /* decoder_pack-p.vhd:199:23  */
  assign n1389_o = n1386_o | n1388_o;
  /* decoder_pack-p.vhd:204:7  */
  assign n1391_o = opc_opcode_q == 8'b00010111;
  /* decoder_pack-p.vhd:204:23  */
  assign n1393_o = opc_opcode_q == 8'b00011000;
  /* decoder_pack-p.vhd:204:23  */
  assign n1394_o = n1391_o | n1393_o;
  /* decoder_pack-p.vhd:205:23  */
  assign n1396_o = opc_opcode_q == 8'b00011001;
  /* decoder_pack-p.vhd:205:23  */
  assign n1397_o = n1394_o | n1396_o;
  /* decoder_pack-p.vhd:205:36  */
  assign n1399_o = opc_opcode_q == 8'b00011010;
  /* decoder_pack-p.vhd:205:36  */
  assign n1400_o = n1397_o | n1399_o;
  /* decoder_pack-p.vhd:205:49  */
  assign n1402_o = opc_opcode_q == 8'b00011011;
  /* decoder_pack-p.vhd:205:49  */
  assign n1403_o = n1400_o | n1402_o;
  /* decoder_pack-p.vhd:205:62  */
  assign n1405_o = opc_opcode_q == 8'b00011100;
  /* decoder_pack-p.vhd:205:62  */
  assign n1406_o = n1403_o | n1405_o;
  /* decoder_pack-p.vhd:206:23  */
  assign n1408_o = opc_opcode_q == 8'b00011101;
  /* decoder_pack-p.vhd:206:23  */
  assign n1409_o = n1406_o | n1408_o;
  /* decoder_pack-p.vhd:206:36  */
  assign n1411_o = opc_opcode_q == 8'b00011110;
  /* decoder_pack-p.vhd:206:36  */
  assign n1412_o = n1409_o | n1411_o;
  /* decoder_pack-p.vhd:206:49  */
  assign n1414_o = opc_opcode_q == 8'b00011111;
  /* decoder_pack-p.vhd:206:49  */
  assign n1415_o = n1412_o | n1414_o;
  /* decoder_pack-p.vhd:206:62  */
  assign n1417_o = opc_opcode_q == 8'b00010000;
  /* decoder_pack-p.vhd:206:62  */
  assign n1418_o = n1415_o | n1417_o;
  /* decoder_pack-p.vhd:207:23  */
  assign n1420_o = opc_opcode_q == 8'b00010001;
  /* decoder_pack-p.vhd:207:23  */
  assign n1421_o = n1418_o | n1420_o;
  /* decoder_pack-p.vhd:211:7  */
  assign n1423_o = opc_opcode_q == 8'b00001000;
  /* decoder_pack-p.vhd:216:7  */
  assign n1425_o = opc_opcode_q == 8'b00010010;
  /* decoder_pack-p.vhd:216:23  */
  assign n1427_o = opc_opcode_q == 8'b00110010;
  /* decoder_pack-p.vhd:216:23  */
  assign n1428_o = n1425_o | n1427_o;
  /* decoder_pack-p.vhd:216:36  */
  assign n1430_o = opc_opcode_q == 8'b01010010;
  /* decoder_pack-p.vhd:216:36  */
  assign n1431_o = n1428_o | n1430_o;
  /* decoder_pack-p.vhd:216:49  */
  assign n1433_o = opc_opcode_q == 8'b01110010;
  /* decoder_pack-p.vhd:216:49  */
  assign n1434_o = n1431_o | n1433_o;
  /* decoder_pack-p.vhd:216:62  */
  assign n1436_o = opc_opcode_q == 8'b10010010;
  /* decoder_pack-p.vhd:216:62  */
  assign n1437_o = n1434_o | n1436_o;
  /* decoder_pack-p.vhd:217:23  */
  assign n1439_o = opc_opcode_q == 8'b10110010;
  /* decoder_pack-p.vhd:217:23  */
  assign n1440_o = n1437_o | n1439_o;
  /* decoder_pack-p.vhd:217:36  */
  assign n1442_o = opc_opcode_q == 8'b11010010;
  /* decoder_pack-p.vhd:217:36  */
  assign n1443_o = n1440_o | n1442_o;
  /* decoder_pack-p.vhd:217:49  */
  assign n1445_o = opc_opcode_q == 8'b11110010;
  /* decoder_pack-p.vhd:217:49  */
  assign n1446_o = n1443_o | n1445_o;
  /* decoder_pack-p.vhd:222:7  */
  assign n1448_o = opc_opcode_q == 8'b11110110;
  /* decoder_pack-p.vhd:222:23  */
  assign n1450_o = opc_opcode_q == 8'b11100110;
  /* decoder_pack-p.vhd:222:23  */
  assign n1451_o = n1448_o | n1450_o;
  /* decoder_pack-p.vhd:228:7  */
  assign n1453_o = opc_opcode_q == 8'b10110110;
  /* decoder_pack-p.vhd:228:23  */
  assign n1455_o = opc_opcode_q == 8'b01110110;
  /* decoder_pack-p.vhd:228:23  */
  assign n1456_o = n1453_o | n1455_o;
  /* decoder_pack-p.vhd:234:7  */
  assign n1458_o = opc_opcode_q == 8'b00000100;
  /* decoder_pack-p.vhd:234:23  */
  assign n1460_o = opc_opcode_q == 8'b00100100;
  /* decoder_pack-p.vhd:234:23  */
  assign n1461_o = n1458_o | n1460_o;
  /* decoder_pack-p.vhd:234:36  */
  assign n1463_o = opc_opcode_q == 8'b01000100;
  /* decoder_pack-p.vhd:234:36  */
  assign n1464_o = n1461_o | n1463_o;
  /* decoder_pack-p.vhd:234:49  */
  assign n1466_o = opc_opcode_q == 8'b01100100;
  /* decoder_pack-p.vhd:234:49  */
  assign n1467_o = n1464_o | n1466_o;
  /* decoder_pack-p.vhd:234:62  */
  assign n1469_o = opc_opcode_q == 8'b10000100;
  /* decoder_pack-p.vhd:234:62  */
  assign n1470_o = n1467_o | n1469_o;
  /* decoder_pack-p.vhd:235:23  */
  assign n1472_o = opc_opcode_q == 8'b10100100;
  /* decoder_pack-p.vhd:235:23  */
  assign n1473_o = n1470_o | n1472_o;
  /* decoder_pack-p.vhd:235:36  */
  assign n1475_o = opc_opcode_q == 8'b11000100;
  /* decoder_pack-p.vhd:235:36  */
  assign n1476_o = n1473_o | n1475_o;
  /* decoder_pack-p.vhd:235:49  */
  assign n1478_o = opc_opcode_q == 8'b11100100;
  /* decoder_pack-p.vhd:235:49  */
  assign n1479_o = n1476_o | n1478_o;
  /* decoder_pack-p.vhd:240:7  */
  assign n1481_o = opc_opcode_q == 8'b10110011;
  /* decoder_pack-p.vhd:245:7  */
  assign n1483_o = opc_opcode_q == 8'b10000110;
  /* decoder_pack-p.vhd:250:7  */
  assign n1485_o = opc_opcode_q == 8'b00100110;
  /* decoder_pack-p.vhd:250:23  */
  assign n1487_o = opc_opcode_q == 8'b01000110;
  /* decoder_pack-p.vhd:250:23  */
  assign n1488_o = n1485_o | n1487_o;
  /* decoder_pack-p.vhd:251:23  */
  assign n1490_o = opc_opcode_q == 8'b00110110;
  /* decoder_pack-p.vhd:251:23  */
  assign n1491_o = n1488_o | n1490_o;
  /* decoder_pack-p.vhd:252:23  */
  assign n1493_o = opc_opcode_q == 8'b01010110;
  /* decoder_pack-p.vhd:252:23  */
  assign n1494_o = n1491_o | n1493_o;
  /* decoder_pack-p.vhd:258:7  */
  assign n1496_o = opc_opcode_q == 8'b00010110;
  /* decoder_pack-p.vhd:263:7  */
  assign n1498_o = opc_opcode_q == 8'b10010110;
  /* decoder_pack-p.vhd:263:23  */
  assign n1500_o = opc_opcode_q == 8'b11000110;
  /* decoder_pack-p.vhd:263:23  */
  assign n1501_o = n1498_o | n1500_o;
  /* decoder_pack-p.vhd:269:7  */
  assign n1503_o = opc_opcode_q == 8'b00100011;
  /* decoder_pack-p.vhd:274:7  */
  assign n1505_o = opc_opcode_q == 8'b11000111;
  /* decoder_pack-p.vhd:278:7  */
  assign n1507_o = opc_opcode_q == 8'b11111000;
  /* decoder_pack-p.vhd:278:23  */
  assign n1509_o = opc_opcode_q == 8'b11111001;
  /* decoder_pack-p.vhd:278:23  */
  assign n1510_o = n1507_o | n1509_o;
  /* decoder_pack-p.vhd:278:36  */
  assign n1512_o = opc_opcode_q == 8'b11111010;
  /* decoder_pack-p.vhd:278:36  */
  assign n1513_o = n1510_o | n1512_o;
  /* decoder_pack-p.vhd:278:49  */
  assign n1515_o = opc_opcode_q == 8'b11111011;
  /* decoder_pack-p.vhd:278:49  */
  assign n1516_o = n1513_o | n1515_o;
  /* decoder_pack-p.vhd:278:62  */
  assign n1518_o = opc_opcode_q == 8'b11111100;
  /* decoder_pack-p.vhd:278:62  */
  assign n1519_o = n1516_o | n1518_o;
  /* decoder_pack-p.vhd:279:23  */
  assign n1521_o = opc_opcode_q == 8'b11111101;
  /* decoder_pack-p.vhd:279:23  */
  assign n1522_o = n1519_o | n1521_o;
  /* decoder_pack-p.vhd:279:36  */
  assign n1524_o = opc_opcode_q == 8'b11111110;
  /* decoder_pack-p.vhd:279:36  */
  assign n1525_o = n1522_o | n1524_o;
  /* decoder_pack-p.vhd:279:49  */
  assign n1527_o = opc_opcode_q == 8'b11111111;
  /* decoder_pack-p.vhd:279:49  */
  assign n1528_o = n1525_o | n1527_o;
  /* decoder_pack-p.vhd:279:62  */
  assign n1530_o = opc_opcode_q == 8'b11110000;
  /* decoder_pack-p.vhd:279:62  */
  assign n1531_o = n1528_o | n1530_o;
  /* decoder_pack-p.vhd:280:23  */
  assign n1533_o = opc_opcode_q == 8'b11110001;
  /* decoder_pack-p.vhd:280:23  */
  assign n1534_o = n1531_o | n1533_o;
  /* decoder_pack-p.vhd:284:7  */
  assign n1536_o = opc_opcode_q == 8'b11010111;
  /* decoder_pack-p.vhd:288:7  */
  assign n1538_o = opc_opcode_q == 8'b10101000;
  /* decoder_pack-p.vhd:288:23  */
  assign n1540_o = opc_opcode_q == 8'b10101001;
  /* decoder_pack-p.vhd:288:23  */
  assign n1541_o = n1538_o | n1540_o;
  /* decoder_pack-p.vhd:288:36  */
  assign n1543_o = opc_opcode_q == 8'b10101010;
  /* decoder_pack-p.vhd:288:36  */
  assign n1544_o = n1541_o | n1543_o;
  /* decoder_pack-p.vhd:288:49  */
  assign n1546_o = opc_opcode_q == 8'b10101011;
  /* decoder_pack-p.vhd:288:49  */
  assign n1547_o = n1544_o | n1546_o;
  /* decoder_pack-p.vhd:288:62  */
  assign n1549_o = opc_opcode_q == 8'b10101100;
  /* decoder_pack-p.vhd:288:62  */
  assign n1550_o = n1547_o | n1549_o;
  /* decoder_pack-p.vhd:289:23  */
  assign n1552_o = opc_opcode_q == 8'b10101101;
  /* decoder_pack-p.vhd:289:23  */
  assign n1553_o = n1550_o | n1552_o;
  /* decoder_pack-p.vhd:289:36  */
  assign n1555_o = opc_opcode_q == 8'b10101110;
  /* decoder_pack-p.vhd:289:36  */
  assign n1556_o = n1553_o | n1555_o;
  /* decoder_pack-p.vhd:289:49  */
  assign n1558_o = opc_opcode_q == 8'b10101111;
  /* decoder_pack-p.vhd:289:49  */
  assign n1559_o = n1556_o | n1558_o;
  /* decoder_pack-p.vhd:289:62  */
  assign n1561_o = opc_opcode_q == 8'b10100000;
  /* decoder_pack-p.vhd:289:62  */
  assign n1562_o = n1559_o | n1561_o;
  /* decoder_pack-p.vhd:290:23  */
  assign n1564_o = opc_opcode_q == 8'b10100001;
  /* decoder_pack-p.vhd:290:23  */
  assign n1565_o = n1562_o | n1564_o;
  /* decoder_pack-p.vhd:294:7  */
  assign n1567_o = opc_opcode_q == 8'b10111000;
  /* decoder_pack-p.vhd:294:23  */
  assign n1569_o = opc_opcode_q == 8'b10111001;
  /* decoder_pack-p.vhd:294:23  */
  assign n1570_o = n1567_o | n1569_o;
  /* decoder_pack-p.vhd:294:36  */
  assign n1572_o = opc_opcode_q == 8'b10111010;
  /* decoder_pack-p.vhd:294:36  */
  assign n1573_o = n1570_o | n1572_o;
  /* decoder_pack-p.vhd:294:49  */
  assign n1575_o = opc_opcode_q == 8'b10111011;
  /* decoder_pack-p.vhd:294:49  */
  assign n1576_o = n1573_o | n1575_o;
  /* decoder_pack-p.vhd:294:62  */
  assign n1578_o = opc_opcode_q == 8'b10111100;
  /* decoder_pack-p.vhd:294:62  */
  assign n1579_o = n1576_o | n1578_o;
  /* decoder_pack-p.vhd:295:23  */
  assign n1581_o = opc_opcode_q == 8'b10111101;
  /* decoder_pack-p.vhd:295:23  */
  assign n1582_o = n1579_o | n1581_o;
  /* decoder_pack-p.vhd:295:36  */
  assign n1584_o = opc_opcode_q == 8'b10111110;
  /* decoder_pack-p.vhd:295:36  */
  assign n1585_o = n1582_o | n1584_o;
  /* decoder_pack-p.vhd:295:49  */
  assign n1587_o = opc_opcode_q == 8'b10111111;
  /* decoder_pack-p.vhd:295:49  */
  assign n1588_o = n1585_o | n1587_o;
  /* decoder_pack-p.vhd:295:62  */
  assign n1590_o = opc_opcode_q == 8'b10110000;
  /* decoder_pack-p.vhd:295:62  */
  assign n1591_o = n1588_o | n1590_o;
  /* decoder_pack-p.vhd:296:23  */
  assign n1593_o = opc_opcode_q == 8'b10110001;
  /* decoder_pack-p.vhd:296:23  */
  assign n1594_o = n1591_o | n1593_o;
  /* decoder_pack-p.vhd:301:7  */
  assign n1596_o = opc_opcode_q == 8'b01100010;
  /* decoder_pack-p.vhd:301:23  */
  assign n1598_o = opc_opcode_q == 8'b01000010;
  /* decoder_pack-p.vhd:301:23  */
  assign n1599_o = n1596_o | n1598_o;
  /* decoder_pack-p.vhd:306:7  */
  assign n1601_o = opc_opcode_q == 8'b00001100;
  /* decoder_pack-p.vhd:306:23  */
  assign n1603_o = opc_opcode_q == 8'b00001101;
  /* decoder_pack-p.vhd:306:23  */
  assign n1604_o = n1601_o | n1603_o;
  /* decoder_pack-p.vhd:306:36  */
  assign n1606_o = opc_opcode_q == 8'b00001110;
  /* decoder_pack-p.vhd:306:36  */
  assign n1607_o = n1604_o | n1606_o;
  /* decoder_pack-p.vhd:306:49  */
  assign n1609_o = opc_opcode_q == 8'b00001111;
  /* decoder_pack-p.vhd:306:49  */
  assign n1610_o = n1607_o | n1609_o;
  /* decoder_pack-p.vhd:311:7  */
  assign n1612_o = opc_opcode_q == 8'b10100011;
  /* decoder_pack-p.vhd:311:23  */
  assign n1614_o = opc_opcode_q == 8'b11100011;
  /* decoder_pack-p.vhd:311:23  */
  assign n1615_o = n1612_o | n1614_o;
  /* decoder_pack-p.vhd:317:7  */
  assign n1617_o = opc_opcode_q == 8'b10000000;
  /* decoder_pack-p.vhd:317:23  */
  assign n1619_o = opc_opcode_q == 8'b10000001;
  /* decoder_pack-p.vhd:317:23  */
  assign n1620_o = n1617_o | n1619_o;
  /* decoder_pack-p.vhd:317:36  */
  assign n1622_o = opc_opcode_q == 8'b10010000;
  /* decoder_pack-p.vhd:317:36  */
  assign n1623_o = n1620_o | n1622_o;
  /* decoder_pack-p.vhd:318:23  */
  assign n1625_o = opc_opcode_q == 8'b10010001;
  /* decoder_pack-p.vhd:318:23  */
  assign n1626_o = n1623_o | n1625_o;
  /* decoder_pack-p.vhd:323:7  */
  assign n1628_o = opc_opcode_q == 8'b00000000;
  /* decoder_pack-p.vhd:327:7  */
  assign n1630_o = opc_opcode_q == 8'b01001000;
  /* decoder_pack-p.vhd:327:23  */
  assign n1632_o = opc_opcode_q == 8'b01001001;
  /* decoder_pack-p.vhd:327:23  */
  assign n1633_o = n1630_o | n1632_o;
  /* decoder_pack-p.vhd:327:36  */
  assign n1635_o = opc_opcode_q == 8'b01001010;
  /* decoder_pack-p.vhd:327:36  */
  assign n1636_o = n1633_o | n1635_o;
  /* decoder_pack-p.vhd:327:49  */
  assign n1638_o = opc_opcode_q == 8'b01001011;
  /* decoder_pack-p.vhd:327:49  */
  assign n1639_o = n1636_o | n1638_o;
  /* decoder_pack-p.vhd:327:62  */
  assign n1641_o = opc_opcode_q == 8'b01001100;
  /* decoder_pack-p.vhd:327:62  */
  assign n1642_o = n1639_o | n1641_o;
  /* decoder_pack-p.vhd:328:23  */
  assign n1644_o = opc_opcode_q == 8'b01001101;
  /* decoder_pack-p.vhd:328:23  */
  assign n1645_o = n1642_o | n1644_o;
  /* decoder_pack-p.vhd:328:36  */
  assign n1647_o = opc_opcode_q == 8'b01001110;
  /* decoder_pack-p.vhd:328:36  */
  assign n1648_o = n1645_o | n1647_o;
  /* decoder_pack-p.vhd:328:49  */
  assign n1650_o = opc_opcode_q == 8'b01001111;
  /* decoder_pack-p.vhd:328:49  */
  assign n1651_o = n1648_o | n1650_o;
  /* decoder_pack-p.vhd:328:62  */
  assign n1653_o = opc_opcode_q == 8'b01000000;
  /* decoder_pack-p.vhd:328:62  */
  assign n1654_o = n1651_o | n1653_o;
  /* decoder_pack-p.vhd:329:23  */
  assign n1656_o = opc_opcode_q == 8'b01000001;
  /* decoder_pack-p.vhd:329:23  */
  assign n1657_o = n1654_o | n1656_o;
  /* decoder_pack-p.vhd:333:7  */
  assign n1659_o = opc_opcode_q == 8'b01000011;
  /* decoder_pack-p.vhd:338:7  */
  assign n1661_o = opc_opcode_q == 8'b10001000;
  /* decoder_pack-p.vhd:338:23  */
  assign n1663_o = opc_opcode_q == 8'b10001001;
  /* decoder_pack-p.vhd:338:23  */
  assign n1664_o = n1661_o | n1663_o;
  /* decoder_pack-p.vhd:339:23  */
  assign n1666_o = opc_opcode_q == 8'b10001010;
  /* decoder_pack-p.vhd:339:23  */
  assign n1667_o = n1664_o | n1666_o;
  /* decoder_pack-p.vhd:344:7  */
  assign n1669_o = opc_opcode_q == 8'b00111100;
  /* decoder_pack-p.vhd:344:23  */
  assign n1671_o = opc_opcode_q == 8'b00111101;
  /* decoder_pack-p.vhd:344:23  */
  assign n1672_o = n1669_o | n1671_o;
  /* decoder_pack-p.vhd:344:36  */
  assign n1674_o = opc_opcode_q == 8'b00111110;
  /* decoder_pack-p.vhd:344:36  */
  assign n1675_o = n1672_o | n1674_o;
  /* decoder_pack-p.vhd:344:49  */
  assign n1677_o = opc_opcode_q == 8'b00111111;
  /* decoder_pack-p.vhd:344:49  */
  assign n1678_o = n1675_o | n1677_o;
  /* decoder_pack-p.vhd:344:62  */
  assign n1680_o = opc_opcode_q == 8'b10011100;
  /* decoder_pack-p.vhd:344:62  */
  assign n1681_o = n1678_o | n1680_o;
  /* decoder_pack-p.vhd:345:23  */
  assign n1683_o = opc_opcode_q == 8'b10011101;
  /* decoder_pack-p.vhd:345:23  */
  assign n1684_o = n1681_o | n1683_o;
  /* decoder_pack-p.vhd:345:36  */
  assign n1686_o = opc_opcode_q == 8'b10011110;
  /* decoder_pack-p.vhd:345:36  */
  assign n1687_o = n1684_o | n1686_o;
  /* decoder_pack-p.vhd:345:49  */
  assign n1689_o = opc_opcode_q == 8'b10011111;
  /* decoder_pack-p.vhd:345:49  */
  assign n1690_o = n1687_o | n1689_o;
  /* decoder_pack-p.vhd:345:62  */
  assign n1692_o = opc_opcode_q == 8'b10001100;
  /* decoder_pack-p.vhd:345:62  */
  assign n1693_o = n1690_o | n1692_o;
  /* decoder_pack-p.vhd:346:23  */
  assign n1695_o = opc_opcode_q == 8'b10001101;
  /* decoder_pack-p.vhd:346:23  */
  assign n1696_o = n1693_o | n1695_o;
  /* decoder_pack-p.vhd:346:36  */
  assign n1698_o = opc_opcode_q == 8'b10001110;
  /* decoder_pack-p.vhd:346:36  */
  assign n1699_o = n1696_o | n1698_o;
  /* decoder_pack-p.vhd:346:49  */
  assign n1701_o = opc_opcode_q == 8'b10001111;
  /* decoder_pack-p.vhd:346:49  */
  assign n1702_o = n1699_o | n1701_o;
  /* decoder_pack-p.vhd:351:7  */
  assign n1704_o = opc_opcode_q == 8'b00111001;
  /* decoder_pack-p.vhd:351:23  */
  assign n1706_o = opc_opcode_q == 8'b00111010;
  /* decoder_pack-p.vhd:351:23  */
  assign n1707_o = n1704_o | n1706_o;
  /* decoder_pack-p.vhd:351:36  */
  assign n1709_o = opc_opcode_q == 8'b00000010;
  /* decoder_pack-p.vhd:351:36  */
  assign n1710_o = n1707_o | n1709_o;
  /* decoder_pack-p.vhd:357:7  */
  assign n1712_o = opc_opcode_q == 8'b10000011;
  /* decoder_pack-p.vhd:357:23  */
  assign n1714_o = opc_opcode_q == 8'b10010011;
  /* decoder_pack-p.vhd:357:23  */
  assign n1715_o = n1712_o | n1714_o;
  /* decoder_pack-p.vhd:363:7  */
  assign n1717_o = opc_opcode_q == 8'b11100111;
  /* decoder_pack-p.vhd:363:23  */
  assign n1719_o = opc_opcode_q == 8'b11110111;
  /* decoder_pack-p.vhd:363:23  */
  assign n1720_o = n1717_o | n1719_o;
  /* decoder_pack-p.vhd:368:7  */
  assign n1722_o = opc_opcode_q == 8'b01110111;
  /* decoder_pack-p.vhd:368:23  */
  assign n1724_o = opc_opcode_q == 8'b01100111;
  /* decoder_pack-p.vhd:368:23  */
  assign n1725_o = n1722_o | n1724_o;
  /* decoder_pack-p.vhd:373:7  */
  assign n1727_o = opc_opcode_q == 8'b11100101;
  /* decoder_pack-p.vhd:373:23  */
  assign n1729_o = opc_opcode_q == 8'b11110101;
  /* decoder_pack-p.vhd:373:23  */
  assign n1730_o = n1727_o | n1729_o;
  /* decoder_pack-p.vhd:378:7  */
  assign n1732_o = opc_opcode_q == 8'b11000101;
  /* decoder_pack-p.vhd:378:23  */
  assign n1734_o = opc_opcode_q == 8'b11010101;
  /* decoder_pack-p.vhd:378:23  */
  assign n1735_o = n1732_o | n1734_o;
  /* decoder_pack-p.vhd:383:7  */
  assign n1737_o = opc_opcode_q == 8'b01100101;
  /* decoder_pack-p.vhd:387:7  */
  assign n1739_o = opc_opcode_q == 8'b01000101;
  /* decoder_pack-p.vhd:387:23  */
  assign n1741_o = opc_opcode_q == 8'b01010101;
  /* decoder_pack-p.vhd:387:23  */
  assign n1742_o = n1739_o | n1741_o;
  /* decoder_pack-p.vhd:392:7  */
  assign n1744_o = opc_opcode_q == 8'b01000111;
  /* decoder_pack-p.vhd:396:7  */
  assign n1746_o = opc_opcode_q == 8'b00101000;
  /* decoder_pack-p.vhd:396:23  */
  assign n1748_o = opc_opcode_q == 8'b00101001;
  /* decoder_pack-p.vhd:396:23  */
  assign n1749_o = n1746_o | n1748_o;
  /* decoder_pack-p.vhd:396:36  */
  assign n1751_o = opc_opcode_q == 8'b00101010;
  /* decoder_pack-p.vhd:396:36  */
  assign n1752_o = n1749_o | n1751_o;
  /* decoder_pack-p.vhd:396:49  */
  assign n1754_o = opc_opcode_q == 8'b00101011;
  /* decoder_pack-p.vhd:396:49  */
  assign n1755_o = n1752_o | n1754_o;
  /* decoder_pack-p.vhd:396:62  */
  assign n1757_o = opc_opcode_q == 8'b00101100;
  /* decoder_pack-p.vhd:396:62  */
  assign n1758_o = n1755_o | n1757_o;
  /* decoder_pack-p.vhd:397:23  */
  assign n1760_o = opc_opcode_q == 8'b00101101;
  /* decoder_pack-p.vhd:397:23  */
  assign n1761_o = n1758_o | n1760_o;
  /* decoder_pack-p.vhd:397:36  */
  assign n1763_o = opc_opcode_q == 8'b00101110;
  /* decoder_pack-p.vhd:397:36  */
  assign n1764_o = n1761_o | n1763_o;
  /* decoder_pack-p.vhd:397:49  */
  assign n1766_o = opc_opcode_q == 8'b00101111;
  /* decoder_pack-p.vhd:397:49  */
  assign n1767_o = n1764_o | n1766_o;
  /* decoder_pack-p.vhd:397:62  */
  assign n1769_o = opc_opcode_q == 8'b00100000;
  /* decoder_pack-p.vhd:397:62  */
  assign n1770_o = n1767_o | n1769_o;
  /* decoder_pack-p.vhd:398:23  */
  assign n1772_o = opc_opcode_q == 8'b00100001;
  /* decoder_pack-p.vhd:398:23  */
  assign n1773_o = n1770_o | n1772_o;
  /* decoder_pack-p.vhd:398:36  */
  assign n1775_o = opc_opcode_q == 8'b00110000;
  /* decoder_pack-p.vhd:398:36  */
  assign n1776_o = n1773_o | n1775_o;
  /* decoder_pack-p.vhd:399:23  */
  assign n1778_o = opc_opcode_q == 8'b00110001;
  /* decoder_pack-p.vhd:399:23  */
  assign n1779_o = n1776_o | n1778_o;
  /* decoder_pack-p.vhd:403:7  */
  assign n1781_o = opc_opcode_q == 8'b11011000;
  /* decoder_pack-p.vhd:403:23  */
  assign n1783_o = opc_opcode_q == 8'b11011001;
  /* decoder_pack-p.vhd:403:23  */
  assign n1784_o = n1781_o | n1783_o;
  /* decoder_pack-p.vhd:403:36  */
  assign n1786_o = opc_opcode_q == 8'b11011010;
  /* decoder_pack-p.vhd:403:36  */
  assign n1787_o = n1784_o | n1786_o;
  /* decoder_pack-p.vhd:403:49  */
  assign n1789_o = opc_opcode_q == 8'b11011011;
  /* decoder_pack-p.vhd:403:49  */
  assign n1790_o = n1787_o | n1789_o;
  /* decoder_pack-p.vhd:403:62  */
  assign n1792_o = opc_opcode_q == 8'b11011100;
  /* decoder_pack-p.vhd:403:62  */
  assign n1793_o = n1790_o | n1792_o;
  /* decoder_pack-p.vhd:404:23  */
  assign n1795_o = opc_opcode_q == 8'b11011101;
  /* decoder_pack-p.vhd:404:23  */
  assign n1796_o = n1793_o | n1795_o;
  /* decoder_pack-p.vhd:404:36  */
  assign n1798_o = opc_opcode_q == 8'b11011110;
  /* decoder_pack-p.vhd:404:36  */
  assign n1799_o = n1796_o | n1798_o;
  /* decoder_pack-p.vhd:404:49  */
  assign n1801_o = opc_opcode_q == 8'b11011111;
  /* decoder_pack-p.vhd:404:49  */
  assign n1802_o = n1799_o | n1801_o;
  /* decoder_pack-p.vhd:404:62  */
  assign n1804_o = opc_opcode_q == 8'b11010000;
  /* decoder_pack-p.vhd:404:62  */
  assign n1805_o = n1802_o | n1804_o;
  /* decoder_pack-p.vhd:405:23  */
  assign n1807_o = opc_opcode_q == 8'b11010001;
  /* decoder_pack-p.vhd:405:23  */
  assign n1808_o = n1805_o | n1807_o;
  /* decoder_pack-p.vhd:409:7  */
  assign n1810_o = opc_opcode_q == 8'b11010011;
  assign n1811_o = {n1810_o, n1808_o, n1779_o, n1744_o, n1742_o, n1737_o, n1735_o, n1730_o, n1725_o, n1720_o, n1715_o, n1710_o, n1702_o, n1667_o, n1659_o, n1657_o, n1628_o, n1626_o, n1615_o, n1610_o, n1599_o, n1594_o, n1565_o, n1536_o, n1534_o, n1505_o, n1503_o, n1501_o, n1496_o, n1494_o, n1483_o, n1481_o, n1479_o, n1456_o, n1451_o, n1446_o, n1423_o, n1421_o, n1389_o, n1384_o, n1382_o, n1359_o, n1354_o, n1349_o, n1323_o, n1321_o, n1316_o, n1314_o, n1312_o, n1307_o, n1305_o, n1303_o, n1280_o, n1272_o, n1270_o, n1241_o, n1236_o};
  /* decoder_pack-p.vhd:103:5  */
  always @*
    case (n1811_o)
      57'b100000000000000000000000000000000000000000000000000000000: n1870_o = 6'b111000;
      57'b010000000000000000000000000000000000000000000000000000000: n1870_o = 6'b110111;
      57'b001000000000000000000000000000000000000000000000000000000: n1870_o = 6'b110110;
      57'b000100000000000000000000000000000000000000000000000000000: n1870_o = 6'b110101;
      57'b000010000000000000000000000000000000000000000000000000000: n1870_o = 6'b110100;
      57'b000001000000000000000000000000000000000000000000000000000: n1870_o = 6'b110011;
      57'b000000100000000000000000000000000000000000000000000000000: n1870_o = 6'b110010;
      57'b000000010000000000000000000000000000000000000000000000000: n1870_o = 6'b110001;
      57'b000000001000000000000000000000000000000000000000000000000: n1870_o = 6'b110000;
      57'b000000000100000000000000000000000000000000000000000000000: n1870_o = 6'b101111;
      57'b000000000010000000000000000000000000000000000000000000000: n1870_o = 6'b101110;
      57'b000000000001000000000000000000000000000000000000000000000: n1870_o = 6'b101101;
      57'b000000000000100000000000000000000000000000000000000000000: n1870_o = 6'b101100;
      57'b000000000000010000000000000000000000000000000000000000000: n1870_o = 6'b101011;
      57'b000000000000001000000000000000000000000000000000000000000: n1870_o = 6'b101010;
      57'b000000000000000100000000000000000000000000000000000000000: n1870_o = 6'b101001;
      57'b000000000000000010000000000000000000000000000000000000000: n1870_o = 6'b101000;
      57'b000000000000000001000000000000000000000000000000000000000: n1870_o = 6'b100111;
      57'b000000000000000000100000000000000000000000000000000000000: n1870_o = 6'b100110;
      57'b000000000000000000010000000000000000000000000000000000000: n1870_o = 6'b100101;
      57'b000000000000000000001000000000000000000000000000000000000: n1870_o = 6'b100100;
      57'b000000000000000000000100000000000000000000000000000000000: n1870_o = 6'b100011;
      57'b000000000000000000000010000000000000000000000000000000000: n1870_o = 6'b100010;
      57'b000000000000000000000001000000000000000000000000000000000: n1870_o = 6'b100001;
      57'b000000000000000000000000100000000000000000000000000000000: n1870_o = 6'b100000;
      57'b000000000000000000000000010000000000000000000000000000000: n1870_o = 6'b011111;
      57'b000000000000000000000000001000000000000000000000000000000: n1870_o = 6'b011110;
      57'b000000000000000000000000000100000000000000000000000000000: n1870_o = 6'b011101;
      57'b000000000000000000000000000010000000000000000000000000000: n1870_o = 6'b011100;
      57'b000000000000000000000000000001000000000000000000000000000: n1870_o = 6'b011011;
      57'b000000000000000000000000000000100000000000000000000000000: n1870_o = 6'b011010;
      57'b000000000000000000000000000000010000000000000000000000000: n1870_o = 6'b011001;
      57'b000000000000000000000000000000001000000000000000000000000: n1870_o = 6'b011000;
      57'b000000000000000000000000000000000100000000000000000000000: n1870_o = 6'b010111;
      57'b000000000000000000000000000000000010000000000000000000000: n1870_o = 6'b010110;
      57'b000000000000000000000000000000000001000000000000000000000: n1870_o = 6'b010101;
      57'b000000000000000000000000000000000000100000000000000000000: n1870_o = 6'b010100;
      57'b000000000000000000000000000000000000010000000000000000000: n1870_o = 6'b010011;
      57'b000000000000000000000000000000000000001000000000000000000: n1870_o = 6'b010010;
      57'b000000000000000000000000000000000000000100000000000000000: n1870_o = 6'b010001;
      57'b000000000000000000000000000000000000000010000000000000000: n1870_o = 6'b010000;
      57'b000000000000000000000000000000000000000001000000000000000: n1870_o = 6'b001111;
      57'b000000000000000000000000000000000000000000100000000000000: n1870_o = 6'b001110;
      57'b000000000000000000000000000000000000000000010000000000000: n1870_o = 6'b001101;
      57'b000000000000000000000000000000000000000000001000000000000: n1870_o = 6'b001100;
      57'b000000000000000000000000000000000000000000000100000000000: n1870_o = 6'b001011;
      57'b000000000000000000000000000000000000000000000010000000000: n1870_o = 6'b001010;
      57'b000000000000000000000000000000000000000000000001000000000: n1870_o = 6'b001001;
      57'b000000000000000000000000000000000000000000000000100000000: n1870_o = 6'b001000;
      57'b000000000000000000000000000000000000000000000000010000000: n1870_o = 6'b000111;
      57'b000000000000000000000000000000000000000000000000001000000: n1870_o = 6'b000110;
      57'b000000000000000000000000000000000000000000000000000100000: n1870_o = 6'b000101;
      57'b000000000000000000000000000000000000000000000000000010000: n1870_o = 6'b000100;
      57'b000000000000000000000000000000000000000000000000000001000: n1870_o = 6'b000011;
      57'b000000000000000000000000000000000000000000000000000000100: n1870_o = 6'b000010;
      57'b000000000000000000000000000000000000000000000000000000010: n1870_o = 6'b000001;
      57'b000000000000000000000000000000000000000000000000000000001: n1870_o = 6'b000000;
      default: n1870_o = 6'b101000;
    endcase
  /* decoder_pack-p.vhd:103:5  */
  always @*
    case (n1811_o)
      57'b100000000000000000000000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b010000000000000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000001000000000000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000100000000000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000010000000000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000001000000000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000100000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000100000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000010000000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000001000000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000010000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000100000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000010000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000001000000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000100000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000010000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000001000000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000100000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000010000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000001000000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000000100000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000000010000000000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000000000100000000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000000000001000000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000000000000000000000010000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000000000000000000000001000: n1900_o = 1'b1;
      57'b000000000000000000000000000000000000000000000000000000100: n1900_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n1900_o = 1'b1;
      57'b000000000000000000000000000000000000000000000000000000001: n1900_o = 1'b0;
      default: n1900_o = 1'b0;
    endcase
  assign n1904_o = {n1900_o, n1870_o};
  /* decoder.vhd:276:14  */
  assign n1906_o = ~res_i;
  /* decoder.vhd:288:40  */
  assign n1908_o = mnemonic_rec_s[5:0];
  /* decoder.vhd:285:9  */
  assign n1910_o = opc_inj_int_s ? 8'b00010100 : opc_opcode_q;
  /* decoder.vhd:285:9  */
  assign n1911_o = opc_inj_int_s ? mnemonic_q : n1908_o;
  /* decoder.vhd:283:9  */
  assign n1912_o = opc_read_bus_s ? data_i : n1910_o;
  /* decoder.vhd:283:9  */
  assign n1913_o = opc_read_bus_s ? mnemonic_q : n1911_o;
  /* decoder.vhd:297:39  */
  assign n1923_o = mnemonic_rec_s[6];
  /* decoder.vhd:299:24  */
  assign n1925_o = 1'b1 ? mnemonic_q : n1926_o;
  /* decoder.vhd:300:41  */
  assign n1926_o = mnemonic_rec_s[5:0];
  /* decoder.vhd:318:28  */
  assign int_b_n1927 = int_b_tf_o; // (signal)
  /* decoder.vhd:327:28  */
  assign int_b_n1929 = int_b_tim_int_o; // (signal)
  /* decoder.vhd:330:28  */
  assign int_b_n1930 = int_b_int_pending_o; // (signal)
  /* decoder.vhd:331:28  */
  assign int_b_n1931 = int_b_int_in_progress_o; // (signal)
  /* decoder.vhd:308:3  */
  t48_int int_b (
    .clk_i(clk_i),
    .res_i(res_i),
    .en_clk_i(en_clk_i),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_i),
    .clk_mstate_i(clk_mstate_i),
    .jtf_executed_i(jtf_executed_s),
    .tim_overflow_i(tim_overflow_i),
    .en_tcnti_i(en_tcnti_s),
    .dis_tcnti_i(dis_tcnti_s),
    .int_n_i(int_n_i),
    .ale_i(ale_i),
    .last_cycle_i(last_cycle_s),
    .en_i_i(en_i_s),
    .dis_i_i(dis_i_s),
    .retr_executed_i(retr_executed_s),
    .int_executed_i(int_executed_s),
    .tf_o(int_b_tf_o),
    .ext_int_o(),
    .tim_int_o(int_b_tim_int_o),
    .int_pending_o(int_b_int_pending_o),
    .int_in_progress_o(int_b_int_in_progress_o));
  /* decoder.vhd:334:19  */
  assign n1941_o = ~opc_multi_cycle_s;
  /* decoder.vhd:335:38  */
  assign n1942_o = clk_second_cycle_i & opc_multi_cycle_s;
  /* decoder.vhd:334:41  */
  assign n1943_o = n1941_o | n1942_o;
  /* decoder.vhd:368:26  */
  assign n1946_o = ~clk_second_cycle_i;
  /* decoder.vhd:369:46  */
  assign n1947_o = assert_psen_s & clk_second_cycle_i;
  /* decoder.vhd:368:49  */
  assign n1948_o = n1946_o | n1947_o;
  /* decoder.vhd:374:19  */
  assign n1949_o = ~ea_i;
  /* decoder.vhd:375:16  */
  assign n1950_o = ~int_pending_s;
  /* decoder.vhd:375:13  */
  assign n1953_o = n1950_o ? 1'b1 : 1'b0;
  /* decoder.vhd:380:16  */
  assign n1954_o = ~int_pending_s;
  /* decoder.vhd:380:13  */
  assign n1957_o = n1954_o ? 1'b1 : 1'b0;
  /* decoder.vhd:374:11  */
  assign n1959_o = n1949_o ? n1953_o : 1'b0;
  /* decoder.vhd:374:11  */
  assign n1962_o = n1949_o ? 1'b0 : 1'b1;
  /* decoder.vhd:374:11  */
  assign n1964_o = n1949_o ? 1'b0 : n1957_o;
  /* decoder.vhd:373:9  */
  assign n1966_o = n1948_o ? n1959_o : 1'b0;
  /* decoder.vhd:373:9  */
  assign n1968_o = n1948_o ? n1962_o : 1'b0;
  /* decoder.vhd:373:9  */
  assign n1970_o = n1948_o ? n1964_o : 1'b0;
  /* decoder.vhd:388:12  */
  assign n1971_o = ~clk_second_cycle_i;
  /* decoder.vhd:389:14  */
  assign n1972_o = ~int_pending_s;
  /* decoder.vhd:389:11  */
  assign n1975_o = n1972_o ? 1'b1 : 1'b0;
  /* decoder.vhd:389:11  */
  assign n1978_o = n1972_o ? 1'b0 : 1'b1;
  /* decoder.vhd:388:9  */
  assign n1980_o = n1971_o ? n1975_o : 1'b0;
  /* decoder.vhd:388:9  */
  assign n1982_o = n1971_o ? n1978_o : 1'b0;
  /* decoder.vhd:372:7  */
  assign n1984_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:397:31  */
  assign n1985_o = ~branch_taken_q;
  /* decoder.vhd:397:27  */
  assign n1986_o = n1985_o & n1948_o;
  /* decoder.vhd:398:12  */
  assign n1987_o = ~int_pending_s;
  /* decoder.vhd:397:50  */
  assign n1988_o = n1987_o & n1986_o;
  /* decoder.vhd:397:9  */
  assign n1991_o = n1988_o ? 1'b1 : 1'b0;
  /* decoder.vhd:396:7  */
  assign n1993_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:403:9  */
  assign n1996_o = n1948_o ? 1'b1 : 1'b0;
  /* decoder.vhd:402:7  */
  assign n1998_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:416:14  */
  assign n1999_o = ~clk_second_cycle_i;
  /* decoder.vhd:416:37  */
  assign n2000_o = assert_psen_s & n1999_o;
  /* decoder.vhd:417:13  */
  assign n2001_o = n2000_o | last_cycle_s;
  /* decoder.vhd:415:23  */
  assign n2002_o = n2001_o & ea_i;
  /* decoder.vhd:415:9  */
  assign n2005_o = n2002_o ? 1'b1 : 1'b0;
  /* decoder.vhd:415:9  */
  assign n2008_o = n2002_o ? 1'b1 : 1'b0;
  /* decoder.vhd:415:9  */
  assign n2011_o = n2002_o ? 1'b1 : 1'b0;
  /* decoder.vhd:414:7  */
  assign n2013_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:425:28  */
  assign n2014_o = n1948_o | last_cycle_s;
  /* decoder.vhd:424:23  */
  assign n2015_o = n2014_o & ea_i;
  /* decoder.vhd:428:12  */
  assign n2016_o = ~p2_output_exp_s;
  /* decoder.vhd:425:45  */
  assign n2017_o = n2016_o & n2015_o;
  /* decoder.vhd:430:12  */
  assign n2018_o = ~movx_first_cycle_s;
  /* decoder.vhd:428:32  */
  assign n2019_o = n2018_o & n2017_o;
  /* decoder.vhd:424:9  */
  assign n2022_o = n2019_o ? 1'b1 : 1'b0;
  /* decoder.vhd:423:7  */
  assign n2024_o = clk_mstate_i == 3'b100;
  assign n2025_o = {n2024_o, n2013_o, n1998_o, n1993_o, n1984_o};
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2027_o = 1'b0;
      5'b01000: n2027_o = 1'b0;
      5'b00100: n2027_o = 1'b0;
      5'b00010: n2027_o = 1'b0;
      5'b00001: n2027_o = n1966_o;
      default: n2027_o = 1'b0;
    endcase
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2030_o = 1'b0;
      5'b01000: n2030_o = n2005_o;
      5'b00100: n2030_o = 1'b0;
      5'b00010: n2030_o = 1'b0;
      5'b00001: n2030_o = 1'b0;
      default: n2030_o = 1'b0;
    endcase
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2033_o = 1'b0;
      5'b01000: n2033_o = n2008_o;
      5'b00100: n2033_o = 1'b0;
      5'b00010: n2033_o = 1'b0;
      5'b00001: n2033_o = 1'b0;
      default: n2033_o = 1'b0;
    endcase
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2036_o = n2022_o;
      5'b01000: n2036_o = n2011_o;
      5'b00100: n2036_o = 1'b0;
      5'b00010: n2036_o = 1'b0;
      5'b00001: n2036_o = n1968_o;
      default: n2036_o = 1'b0;
    endcase
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2039_o = 1'b0;
      5'b01000: n2039_o = 1'b0;
      5'b00100: n2039_o = 1'b0;
      5'b00010: n2039_o = 1'b0;
      5'b00001: n2039_o = n1980_o;
      default: n2039_o = 1'b0;
    endcase
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2042_o = 1'b0;
      5'b01000: n2042_o = 1'b0;
      5'b00100: n2042_o = 1'b0;
      5'b00010: n2042_o = 1'b0;
      5'b00001: n2042_o = n1982_o;
      default: n2042_o = 1'b0;
    endcase
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2045_o = 1'b0;
      5'b01000: n2045_o = 1'b0;
      5'b00100: n2045_o = 1'b0;
      5'b00010: n2045_o = n1991_o;
      5'b00001: n2045_o = 1'b0;
      default: n2045_o = 1'b0;
    endcase
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2048_o = 1'b0;
      5'b01000: n2048_o = 1'b0;
      5'b00100: n2048_o = n1996_o;
      5'b00010: n2048_o = 1'b0;
      5'b00001: n2048_o = 1'b0;
      default: n2048_o = 1'b0;
    endcase
  /* decoder.vhd:371:5  */
  always @*
    case (n2025_o)
      5'b10000: n2051_o = 1'b0;
      5'b01000: n2051_o = 1'b0;
      5'b00100: n2051_o = 1'b0;
      5'b00010: n2051_o = 1'b0;
      5'b00001: n2051_o = n1970_o;
      default: n2051_o = 1'b0;
    endcase
  /* decoder.vhd:586:5  */
  assign n2058_o = int_in_progress_s ? 1'b0 : mb_q;
  /* decoder.vhd:593:8  */
  assign n2059_o = ~clk_second_cycle_i;
  /* decoder.vhd:593:48  */
  assign n2061_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:593:31  */
  assign n2062_o = n2061_o & n2059_o;
  /* decoder.vhd:595:22  */
  assign n2063_o = opc_opcode_q[3];
  /* decoder.vhd:596:43  */
  assign n2064_o = opc_opcode_q[2:0];
  /* decoder.vhd:598:50  */
  assign n2065_o = opc_opcode_q[0];
  /* decoder.vhd:598:36  */
  assign n2067_o = {2'b00, n2065_o};
  /* decoder.vhd:595:7  */
  assign n2068_o = n2063_o ? n2064_o : n2067_o;
  assign n2070_o = n2069_o[7:3];
  /* decoder.vhd:593:5  */
  assign n2073_o = n2062_o ? 1'b1 : 1'b0;
  assign n2075_o = {n2070_o, n2068_o};
  /* decoder.vhd:593:5  */
  assign n2077_o = n2062_o ? n2075_o : 8'bX;
  /* decoder.vhd:593:5  */
  assign n2081_o = n2062_o ? 1'b1 : 1'b0;
  /* decoder.vhd:614:28  */
  assign n2083_o = opc_opcode_q[3];
  /* decoder.vhd:614:32  */
  assign n2084_o = ~n2083_o;
  /* decoder.vhd:613:44  */
  assign n2086_o = 1'b0 | n2084_o;
  /* decoder.vhd:613:13  */
  assign n2093_o = n2086_o ? 1'b1 : n2073_o;
  /* decoder.vhd:613:13  */
  assign n2096_o = n2086_o ? 1'b1 : 1'b0;
  /* decoder.vhd:613:13  */
  assign n2099_o = n2086_o ? 2'b00 : 2'b01;
  /* decoder.vhd:612:11  */
  assign n2101_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:619:11  */
  assign n2106_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:626:28  */
  assign n2110_o = opc_opcode_q[4];
  /* decoder.vhd:626:13  */
  assign n2113_o = n2110_o ? 1'b1 : 1'b0;
  /* decoder.vhd:623:11  */
  assign n2115_o = clk_mstate_i == 3'b100;
  assign n2116_o = {n2115_o, n2106_o, n2101_o};
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2119_o = 1'b1;
      3'b010: n2119_o = 1'b0;
      3'b001: n2119_o = 1'b0;
      default: n2119_o = 1'b0;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2122_o = 1'b0;
      3'b010: n2122_o = 1'b1;
      3'b001: n2122_o = 1'b0;
      default: n2122_o = 1'b0;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2125_o = 1'b1;
      3'b010: n2125_o = 1'b0;
      3'b001: n2125_o = 1'b0;
      default: n2125_o = 1'b0;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2126_o = n2073_o;
      3'b010: n2126_o = n2073_o;
      3'b001: n2126_o = n2093_o;
      default: n2126_o = n2073_o;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2129_o = 1'b0;
      3'b010: n2129_o = 1'b1;
      3'b001: n2129_o = n2096_o;
      default: n2129_o = 1'b0;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2132_o = 4'b1010;
      3'b010: n2132_o = 4'b1100;
      3'b001: n2132_o = 4'b1100;
      default: n2132_o = 4'b1100;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2134_o = n2113_o;
      3'b010: n2134_o = 1'b0;
      3'b001: n2134_o = 1'b0;
      default: n2134_o = 1'b0;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2136_o = 2'b01;
      3'b010: n2136_o = 2'b01;
      3'b001: n2136_o = n2099_o;
      default: n2136_o = 2'b01;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2138_o = alu_carry_i;
      3'b010: n2138_o = 1'b0;
      3'b001: n2138_o = 1'b0;
      default: n2138_o = 1'b0;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2141_o = 1'b1;
      3'b010: n2141_o = 1'b0;
      3'b001: n2141_o = 1'b0;
      default: n2141_o = 1'b0;
    endcase
  /* decoder.vhd:610:9  */
  always @*
    case (n2116_o)
      3'b100: n2144_o = 1'b1;
      3'b010: n2144_o = 1'b0;
      3'b001: n2144_o = 1'b0;
      default: n2144_o = 1'b0;
    endcase
  /* decoder.vhd:609:7  */
  assign n2146_o = opc_mnemonic_s == 6'b000000;
  /* decoder.vhd:646:13  */
  assign n2148_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:653:30  */
  assign n2152_o = opc_opcode_q[4];
  /* decoder.vhd:653:15  */
  assign n2155_o = n2152_o ? 1'b1 : 1'b0;
  /* decoder.vhd:650:13  */
  assign n2157_o = clk_mstate_i == 3'b010;
  assign n2158_o = {n2157_o, n2148_o};
  /* decoder.vhd:644:11  */
  always @*
    case (n2158_o)
      2'b10: n2161_o = 1'b1;
      2'b01: n2161_o = 1'b0;
      default: n2161_o = 1'b0;
    endcase
  /* decoder.vhd:644:11  */
  always @*
    case (n2158_o)
      2'b10: n2164_o = 1'b0;
      2'b01: n2164_o = 1'b1;
      default: n2164_o = 1'b0;
    endcase
  /* decoder.vhd:644:11  */
  always @*
    case (n2158_o)
      2'b10: n2167_o = 1'b1;
      2'b01: n2167_o = 1'b0;
      default: n2167_o = 1'b0;
    endcase
  /* decoder.vhd:644:11  */
  always @*
    case (n2158_o)
      2'b10: n2170_o = 4'b1010;
      2'b01: n2170_o = 4'b1100;
      default: n2170_o = 4'b1100;
    endcase
  /* decoder.vhd:644:11  */
  always @*
    case (n2158_o)
      2'b10: n2172_o = n2155_o;
      2'b01: n2172_o = 1'b0;
      default: n2172_o = 1'b0;
    endcase
  /* decoder.vhd:644:11  */
  always @*
    case (n2158_o)
      2'b10: n2174_o = alu_carry_i;
      2'b01: n2174_o = 1'b0;
      default: n2174_o = 1'b0;
    endcase
  /* decoder.vhd:644:11  */
  always @*
    case (n2158_o)
      2'b10: n2177_o = 1'b1;
      2'b01: n2177_o = 1'b0;
      default: n2177_o = 1'b0;
    endcase
  /* decoder.vhd:644:11  */
  always @*
    case (n2158_o)
      2'b10: n2180_o = 1'b1;
      2'b01: n2180_o = 1'b0;
      default: n2180_o = 1'b0;
    endcase
  /* decoder.vhd:643:9  */
  assign n2182_o = clk_second_cycle_i ? n2161_o : 1'b0;
  /* decoder.vhd:643:9  */
  assign n2184_o = clk_second_cycle_i ? n2164_o : 1'b0;
  /* decoder.vhd:643:9  */
  assign n2186_o = clk_second_cycle_i ? n2167_o : 1'b0;
  /* decoder.vhd:643:9  */
  assign n2188_o = clk_second_cycle_i ? n2170_o : 4'b1100;
  /* decoder.vhd:643:9  */
  assign n2190_o = clk_second_cycle_i ? n2172_o : 1'b0;
  /* decoder.vhd:643:9  */
  assign n2192_o = clk_second_cycle_i ? n2174_o : 1'b0;
  /* decoder.vhd:643:9  */
  assign n2194_o = clk_second_cycle_i ? n2177_o : 1'b0;
  /* decoder.vhd:643:9  */
  assign n2196_o = clk_second_cycle_i ? n2180_o : 1'b0;
  /* decoder.vhd:640:7  */
  assign n2198_o = opc_mnemonic_s == 6'b000001;
  /* decoder.vhd:674:28  */
  assign n2199_o = opc_opcode_q[3];
  /* decoder.vhd:674:32  */
  assign n2200_o = ~n2199_o;
  /* decoder.vhd:673:44  */
  assign n2202_o = 1'b0 | n2200_o;
  /* decoder.vhd:673:13  */
  assign n2209_o = n2202_o ? 1'b1 : n2073_o;
  /* decoder.vhd:673:13  */
  assign n2212_o = n2202_o ? 1'b1 : 1'b0;
  /* decoder.vhd:673:13  */
  assign n2215_o = n2202_o ? 2'b00 : 2'b01;
  /* decoder.vhd:672:11  */
  assign n2217_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:679:11  */
  assign n2222_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:683:11  */
  assign n2227_o = clk_mstate_i == 3'b100;
  assign n2228_o = {n2227_o, n2222_o, n2217_o};
  /* decoder.vhd:670:9  */
  always @*
    case (n2228_o)
      3'b100: n2231_o = 1'b1;
      3'b010: n2231_o = 1'b0;
      3'b001: n2231_o = 1'b0;
      default: n2231_o = 1'b0;
    endcase
  /* decoder.vhd:670:9  */
  always @*
    case (n2228_o)
      3'b100: n2234_o = 1'b0;
      3'b010: n2234_o = 1'b1;
      3'b001: n2234_o = 1'b0;
      default: n2234_o = 1'b0;
    endcase
  /* decoder.vhd:670:9  */
  always @*
    case (n2228_o)
      3'b100: n2237_o = 1'b1;
      3'b010: n2237_o = 1'b0;
      3'b001: n2237_o = 1'b0;
      default: n2237_o = 1'b0;
    endcase
  /* decoder.vhd:670:9  */
  always @*
    case (n2228_o)
      3'b100: n2238_o = n2073_o;
      3'b010: n2238_o = n2073_o;
      3'b001: n2238_o = n2209_o;
      default: n2238_o = n2073_o;
    endcase
  /* decoder.vhd:670:9  */
  always @*
    case (n2228_o)
      3'b100: n2241_o = 1'b0;
      3'b010: n2241_o = 1'b1;
      3'b001: n2241_o = n2212_o;
      default: n2241_o = 1'b0;
    endcase
  /* decoder.vhd:670:9  */
  always @*
    case (n2228_o)
      3'b100: n2244_o = 4'b0000;
      3'b010: n2244_o = 4'b1100;
      3'b001: n2244_o = 4'b1100;
      default: n2244_o = 4'b1100;
    endcase
  /* decoder.vhd:670:9  */
  always @*
    case (n2228_o)
      3'b100: n2246_o = 2'b01;
      3'b010: n2246_o = 2'b01;
      3'b001: n2246_o = n2215_o;
      default: n2246_o = 2'b01;
    endcase
  /* decoder.vhd:669:7  */
  assign n2248_o = opc_mnemonic_s == 6'b000010;
  /* decoder.vhd:698:13  */
  assign n2250_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:702:13  */
  assign n2255_o = clk_mstate_i == 3'b010;
  assign n2256_o = {n2255_o, n2250_o};
  /* decoder.vhd:696:11  */
  always @*
    case (n2256_o)
      2'b10: n2259_o = 1'b1;
      2'b01: n2259_o = 1'b0;
      default: n2259_o = 1'b0;
    endcase
  /* decoder.vhd:696:11  */
  always @*
    case (n2256_o)
      2'b10: n2262_o = 1'b0;
      2'b01: n2262_o = 1'b1;
      default: n2262_o = 1'b0;
    endcase
  /* decoder.vhd:696:11  */
  always @*
    case (n2256_o)
      2'b10: n2265_o = 1'b1;
      2'b01: n2265_o = 1'b0;
      default: n2265_o = 1'b0;
    endcase
  /* decoder.vhd:696:11  */
  always @*
    case (n2256_o)
      2'b10: n2268_o = 4'b0000;
      2'b01: n2268_o = 4'b1100;
      default: n2268_o = 4'b1100;
    endcase
  /* decoder.vhd:695:9  */
  assign n2270_o = clk_second_cycle_i ? n2259_o : 1'b0;
  /* decoder.vhd:695:9  */
  assign n2272_o = clk_second_cycle_i ? n2262_o : 1'b0;
  /* decoder.vhd:695:9  */
  assign n2274_o = clk_second_cycle_i ? n2265_o : 1'b0;
  /* decoder.vhd:695:9  */
  assign n2276_o = clk_second_cycle_i ? n2268_o : 4'b1100;
  /* decoder.vhd:692:7  */
  assign n2278_o = opc_mnemonic_s == 6'b000011;
  /* decoder.vhd:716:12  */
  assign n2279_o = ~clk_second_cycle_i;
  /* decoder.vhd:718:27  */
  assign n2281_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:719:28  */
  assign n2282_o = opc_opcode_q[1:0];
  /* decoder.vhd:719:41  */
  assign n2284_o = n2282_o == 2'b00;
  /* decoder.vhd:721:31  */
  assign n2285_o = opc_opcode_q[1];
  /* decoder.vhd:721:35  */
  assign n2286_o = ~n2285_o;
  /* decoder.vhd:721:13  */
  assign n2289_o = n2286_o ? 1'b1 : 1'b0;
  /* decoder.vhd:721:13  */
  assign n2292_o = n2286_o ? 1'b0 : 1'b1;
  /* decoder.vhd:721:13  */
  assign n2295_o = n2286_o ? 1'b1 : 1'b0;
  /* decoder.vhd:721:13  */
  assign n2298_o = n2286_o ? 1'b0 : 1'b1;
  /* decoder.vhd:719:13  */
  assign n2300_o = n2284_o ? 1'b0 : n2289_o;
  /* decoder.vhd:719:13  */
  assign n2302_o = n2284_o ? 1'b0 : n2292_o;
  /* decoder.vhd:719:13  */
  assign n2304_o = n2284_o ? 1'b0 : n2295_o;
  /* decoder.vhd:719:13  */
  assign n2306_o = n2284_o ? 1'b0 : n2298_o;
  /* decoder.vhd:719:13  */
  assign n2309_o = n2284_o ? 1'b1 : 1'b0;
  /* decoder.vhd:718:11  */
  assign n2312_o = n2281_o ? 1'b1 : 1'b0;
  /* decoder.vhd:718:11  */
  assign n2314_o = n2281_o ? n2300_o : 1'b0;
  /* decoder.vhd:718:11  */
  assign n2316_o = n2281_o ? n2302_o : 1'b0;
  /* decoder.vhd:718:11  */
  assign n2318_o = n2281_o ? n2304_o : 1'b0;
  /* decoder.vhd:718:11  */
  assign n2320_o = n2281_o ? n2306_o : 1'b0;
  /* decoder.vhd:718:11  */
  assign n2322_o = n2281_o ? n2309_o : 1'b0;
  /* decoder.vhd:736:13  */
  assign n2324_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:741:13  */
  assign n2326_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:750:30  */
  assign n2327_o = opc_opcode_q[1:0];
  /* decoder.vhd:750:43  */
  assign n2329_o = n2327_o == 2'b00;
  /* decoder.vhd:752:33  */
  assign n2330_o = opc_opcode_q[1];
  /* decoder.vhd:752:37  */
  assign n2331_o = ~n2330_o;
  /* decoder.vhd:752:15  */
  assign n2334_o = n2331_o ? 1'b1 : 1'b0;
  /* decoder.vhd:752:15  */
  assign n2337_o = n2331_o ? 1'b0 : 1'b1;
  /* decoder.vhd:750:15  */
  assign n2340_o = n2329_o ? 1'b1 : 1'b0;
  /* decoder.vhd:750:15  */
  assign n2342_o = n2329_o ? 1'b0 : n2334_o;
  /* decoder.vhd:750:15  */
  assign n2344_o = n2329_o ? 1'b0 : n2337_o;
  /* decoder.vhd:746:13  */
  assign n2346_o = clk_mstate_i == 3'b010;
  assign n2347_o = {n2346_o, n2326_o, n2324_o};
  /* decoder.vhd:733:11  */
  always @*
    case (n2347_o)
      3'b100: n2351_o = 1'b0;
      3'b010: n2351_o = 1'b1;
      3'b001: n2351_o = 1'b1;
      default: n2351_o = 1'b0;
    endcase
  /* decoder.vhd:733:11  */
  always @*
    case (n2347_o)
      3'b100: n2355_o = 1'b1;
      3'b010: n2355_o = 1'b1;
      3'b001: n2355_o = 1'b0;
      default: n2355_o = 1'b0;
    endcase
  /* decoder.vhd:733:11  */
  always @*
    case (n2347_o)
      3'b100: n2357_o = n2340_o;
      3'b010: n2357_o = 1'b0;
      3'b001: n2357_o = 1'b0;
      default: n2357_o = 1'b0;
    endcase
  /* decoder.vhd:733:11  */
  always @*
    case (n2347_o)
      3'b100: n2359_o = n2342_o;
      3'b010: n2359_o = 1'b0;
      3'b001: n2359_o = 1'b0;
      default: n2359_o = 1'b0;
    endcase
  /* decoder.vhd:733:11  */
  always @*
    case (n2347_o)
      3'b100: n2361_o = n2344_o;
      3'b010: n2361_o = 1'b0;
      3'b001: n2361_o = 1'b0;
      default: n2361_o = 1'b0;
    endcase
  /* decoder.vhd:733:11  */
  always @*
    case (n2347_o)
      3'b100: n2364_o = 4'b0000;
      3'b010: n2364_o = 4'b1100;
      3'b001: n2364_o = 4'b1100;
      default: n2364_o = 4'b1100;
    endcase
  /* decoder.vhd:716:9  */
  assign n2366_o = n2279_o ? 1'b0 : n2351_o;
  /* decoder.vhd:716:9  */
  assign n2368_o = n2279_o ? n2312_o : 1'b0;
  /* decoder.vhd:716:9  */
  assign n2370_o = n2279_o ? 1'b0 : n2355_o;
  /* decoder.vhd:716:9  */
  assign n2372_o = n2279_o ? 1'b0 : n2357_o;
  /* decoder.vhd:716:9  */
  assign n2374_o = n2279_o ? 1'b0 : n2359_o;
  /* decoder.vhd:716:9  */
  assign n2376_o = n2279_o ? n2314_o : 1'b0;
  /* decoder.vhd:716:9  */
  assign n2378_o = n2279_o ? 1'b0 : n2361_o;
  /* decoder.vhd:716:9  */
  assign n2380_o = n2279_o ? n2316_o : 1'b0;
  /* decoder.vhd:716:9  */
  assign n2382_o = n2279_o ? 4'b1100 : n2364_o;
  /* decoder.vhd:716:9  */
  assign n2384_o = n2279_o ? n2318_o : 1'b0;
  /* decoder.vhd:716:9  */
  assign n2386_o = n2279_o ? n2320_o : 1'b0;
  /* decoder.vhd:716:9  */
  assign n2388_o = n2279_o ? n2322_o : 1'b0;
  /* decoder.vhd:713:7  */
  assign n2390_o = opc_mnemonic_s == 6'b000100;
  /* decoder.vhd:769:12  */
  assign n2391_o = ~clk_second_cycle_i;
  /* decoder.vhd:782:18  */
  assign n2392_o = ~int_pending_s;
  /* decoder.vhd:782:15  */
  assign n2395_o = n2392_o ? 1'b1 : 1'b0;
  /* decoder.vhd:773:13  */
  assign n2397_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:787:13  */
  assign n2399_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:793:13  */
  assign n2401_o = clk_mstate_i == 3'b100;
  assign n2402_o = {n2401_o, n2399_o, n2397_o};
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2405_o = 1'b1;
      3'b010: n2405_o = n2073_o;
      3'b001: n2405_o = 1'b1;
      default: n2405_o = n2073_o;
    endcase
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2408_o = 1'b0;
      3'b010: n2408_o = 1'b1;
      3'b001: n2408_o = 1'b0;
      default: n2408_o = 1'b0;
    endcase
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2411_o = 1'b1;
      3'b010: n2411_o = 1'b0;
      3'b001: n2411_o = 1'b0;
      default: n2411_o = 1'b0;
    endcase
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2414_o = 1'b1;
      3'b010: n2414_o = 1'b0;
      3'b001: n2414_o = 1'b0;
      default: n2414_o = 1'b0;
    endcase
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2417_o = 1'b0;
      3'b010: n2417_o = 1'b0;
      3'b001: n2417_o = 1'b1;
      default: n2417_o = 1'b0;
    endcase
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2421_o = 2'b11;
      3'b010: n2421_o = 2'b01;
      3'b001: n2421_o = 2'b10;
      default: n2421_o = 2'b01;
    endcase
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2424_o = 1'b1;
      3'b010: n2424_o = 1'b0;
      3'b001: n2424_o = 1'b0;
      default: n2424_o = 1'b0;
    endcase
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2426_o = 1'b0;
      3'b010: n2426_o = 1'b0;
      3'b001: n2426_o = n2395_o;
      default: n2426_o = 1'b0;
    endcase
  /* decoder.vhd:770:11  */
  always @*
    case (n2402_o)
      3'b100: n2430_o = 1'b1;
      3'b010: n2430_o = 1'b1;
      3'b001: n2430_o = 1'b0;
      default: n2430_o = 1'b0;
    endcase
  assign n2435_o = n2432_o[2];
  /* decoder.vhd:816:17  */
  assign n2436_o = tim_int_s ? 1'b1 : n2435_o;
  assign n2437_o = n2432_o[7:3];
  assign n2438_o = {n2437_o, n2436_o, 2'b11};
  /* decoder.vhd:812:15  */
  assign n2439_o = int_pending_s ? n2438_o : n2077_o;
  /* decoder.vhd:812:15  */
  assign n2441_o = int_pending_s ? 1'b1 : n2081_o;
  /* decoder.vhd:809:13  */
  assign n2443_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:825:18  */
  assign n2444_o = ~int_pending_s;
  /* decoder.vhd:827:46  */
  assign n2446_o = {4'b0000, n2058_o};
  /* decoder.vhd:827:67  */
  assign n2447_o = opc_opcode_q[7:5];
  /* decoder.vhd:827:53  */
  assign n2448_o = {n2446_o, n2447_o};
  /* decoder.vhd:825:15  */
  assign n2450_o = n2444_o ? n2448_o : 8'b00000000;
  /* decoder.vhd:825:15  */
  assign n2453_o = n2444_o ? 1'b0 : 1'b1;
  /* decoder.vhd:822:13  */
  assign n2455_o = clk_mstate_i == 3'b001;
  assign n2456_o = {n2455_o, n2443_o};
  /* decoder.vhd:807:11  */
  always @*
    case (n2456_o)
      2'b10: n2459_o = 1'b0;
      2'b01: n2459_o = 1'b1;
      default: n2459_o = 1'b0;
    endcase
  /* decoder.vhd:807:11  */
  always @*
    case (n2456_o)
      2'b10: n2462_o = 1'b1;
      2'b01: n2462_o = 1'b0;
      default: n2462_o = 1'b0;
    endcase
  /* decoder.vhd:807:11  */
  always @*
    case (n2456_o)
      2'b10: n2465_o = 1'b0;
      2'b01: n2465_o = 1'b1;
      default: n2465_o = 1'b0;
    endcase
  /* decoder.vhd:807:11  */
  always @*
    case (n2456_o)
      2'b10: n2466_o = n2450_o;
      2'b01: n2466_o = n2439_o;
      default: n2466_o = n2077_o;
    endcase
  /* decoder.vhd:807:11  */
  always @*
    case (n2456_o)
      2'b10: n2468_o = 1'b1;
      2'b01: n2468_o = n2441_o;
      default: n2468_o = n2081_o;
    endcase
  /* decoder.vhd:807:11  */
  always @*
    case (n2456_o)
      2'b10: n2470_o = n2453_o;
      2'b01: n2470_o = 1'b0;
      default: n2470_o = 1'b0;
    endcase
  /* decoder.vhd:769:9  */
  assign n2471_o = n2391_o ? n2405_o : n2073_o;
  /* decoder.vhd:769:9  */
  assign n2473_o = n2391_o ? 1'b0 : n2459_o;
  /* decoder.vhd:769:9  */
  assign n2475_o = n2391_o ? n2408_o : 1'b0;
  /* decoder.vhd:769:9  */
  assign n2477_o = n2391_o ? 1'b0 : n2462_o;
  /* decoder.vhd:769:9  */
  assign n2479_o = n2391_o ? n2411_o : 1'b0;
  /* decoder.vhd:769:9  */
  assign n2481_o = n2391_o ? n2414_o : 1'b0;
  /* decoder.vhd:769:9  */
  assign n2483_o = n2391_o ? n2417_o : 1'b0;
  /* decoder.vhd:769:9  */
  assign n2485_o = n2391_o ? n2421_o : 2'b01;
  /* decoder.vhd:769:9  */
  assign n2487_o = n2391_o ? n2424_o : 1'b0;
  /* decoder.vhd:769:9  */
  assign n2489_o = n2391_o ? 1'b0 : n2465_o;
  /* decoder.vhd:769:9  */
  assign n2491_o = n2391_o ? n2426_o : 1'b0;
  /* decoder.vhd:769:9  */
  assign n2492_o = n2391_o ? n2077_o : n2466_o;
  /* decoder.vhd:769:9  */
  assign n2493_o = n2391_o ? n2081_o : n2468_o;
  /* decoder.vhd:769:9  */
  assign n2495_o = n2391_o ? n2430_o : 1'b0;
  /* decoder.vhd:769:9  */
  assign n2497_o = n2391_o ? 1'b0 : n2470_o;
  /* decoder.vhd:766:7  */
  assign n2499_o = opc_mnemonic_s == 6'b000101;
  /* decoder.vhd:844:25  */
  assign n2501_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:844:9  */
  assign n2504_o = n2501_o ? 1'b1 : 1'b0;
  /* decoder.vhd:844:9  */
  assign n2507_o = n2501_o ? 1'b1 : 1'b0;
  /* decoder.vhd:844:9  */
  assign n2510_o = n2501_o ? 4'b0100 : 4'b1100;
  /* decoder.vhd:842:7  */
  assign n2512_o = opc_mnemonic_s == 6'b000110;
  /* decoder.vhd:853:25  */
  assign n2514_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:853:9  */
  assign n2517_o = n2514_o ? 1'b1 : 1'b0;
  /* decoder.vhd:851:7  */
  assign n2519_o = opc_mnemonic_s == 6'b000111;
  /* decoder.vhd:861:25  */
  assign n2521_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:862:26  */
  assign n2522_o = opc_opcode_q[5];
  /* decoder.vhd:862:30  */
  assign n2523_o = ~n2522_o;
  /* decoder.vhd:862:11  */
  assign n2526_o = n2523_o ? 1'b1 : 1'b0;
  /* decoder.vhd:862:11  */
  assign n2529_o = n2523_o ? 1'b0 : 1'b1;
  /* decoder.vhd:861:9  */
  assign n2531_o = n2521_o ? n2526_o : 1'b0;
  /* decoder.vhd:861:9  */
  assign n2533_o = n2521_o ? n2529_o : 1'b0;
  /* decoder.vhd:859:7  */
  assign n2535_o = opc_mnemonic_s == 6'b001000;
  /* decoder.vhd:874:25  */
  assign n2537_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:874:9  */
  assign n2540_o = n2537_o ? 1'b1 : 1'b0;
  /* decoder.vhd:874:9  */
  assign n2543_o = n2537_o ? 1'b1 : 1'b0;
  /* decoder.vhd:874:9  */
  assign n2546_o = n2537_o ? 4'b0011 : 4'b1100;
  /* decoder.vhd:872:7  */
  assign n2548_o = opc_mnemonic_s == 6'b001001;
  /* decoder.vhd:883:25  */
  assign n2550_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:884:33  */
  assign n2551_o = ~psw_carry_i;
  /* decoder.vhd:883:9  */
  assign n2553_o = n2550_o ? n2551_o : 1'b0;
  /* decoder.vhd:883:9  */
  assign n2556_o = n2550_o ? 1'b1 : 1'b0;
  /* decoder.vhd:881:7  */
  assign n2558_o = opc_mnemonic_s == 6'b001010;
  /* decoder.vhd:891:25  */
  assign n2560_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:892:26  */
  assign n2561_o = opc_opcode_q[5];
  /* decoder.vhd:892:30  */
  assign n2562_o = ~n2561_o;
  /* decoder.vhd:893:35  */
  assign n2563_o = ~psw_f0_i;
  /* decoder.vhd:892:11  */
  assign n2565_o = n2562_o ? n2563_o : 1'b0;
  /* decoder.vhd:892:11  */
  assign n2568_o = n2562_o ? 1'b1 : 1'b0;
  /* decoder.vhd:892:11  */
  assign n2571_o = n2562_o ? 1'b0 : 1'b1;
  /* decoder.vhd:891:9  */
  assign n2573_o = n2560_o ? n2565_o : 1'b0;
  /* decoder.vhd:891:9  */
  assign n2575_o = n2560_o ? n2568_o : 1'b0;
  /* decoder.vhd:891:9  */
  assign n2577_o = n2560_o ? n2571_o : 1'b0;
  /* decoder.vhd:889:7  */
  assign n2579_o = opc_mnemonic_s == 6'b001011;
  /* decoder.vhd:907:11  */
  assign n2581_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:913:38  */
  assign n2582_o = psw_aux_carry_i | alu_da_overflow_i;
  /* decoder.vhd:913:13  */
  assign n2585_o = n2582_o ? 1'b1 : 1'b0;
  /* decoder.vhd:913:13  */
  assign n2588_o = n2582_o ? 1'b1 : 1'b0;
  /* decoder.vhd:912:11  */
  assign n2590_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:927:13  */
  assign n2593_o = alu_da_overflow_i ? 4'b1010 : 4'b1100;
  /* decoder.vhd:927:13  */
  assign n2595_o = alu_da_overflow_i ? alu_carry_i : 1'b0;
  /* decoder.vhd:924:11  */
  assign n2597_o = clk_mstate_i == 3'b100;
  assign n2598_o = {n2597_o, n2590_o, n2581_o};
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2601_o = 1'b1;
      3'b010: n2601_o = 1'b0;
      3'b001: n2601_o = 1'b0;
      default: n2601_o = 1'b0;
    endcase
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2603_o = 1'b0;
      3'b010: n2603_o = n2585_o;
      3'b001: n2603_o = 1'b0;
      default: n2603_o = 1'b0;
    endcase
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2606_o = 1'b1;
      3'b010: n2606_o = n2588_o;
      3'b001: n2606_o = 1'b0;
      default: n2606_o = 1'b0;
    endcase
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2608_o = n2593_o;
      3'b010: n2608_o = 4'b1010;
      3'b001: n2608_o = 4'b1010;
      default: n2608_o = 4'b1010;
    endcase
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2612_o = 1'b1;
      3'b010: n2612_o = 1'b0;
      3'b001: n2612_o = 1'b0;
      default: n2612_o = 1'b0;
    endcase
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2615_o = 1'b0;
      3'b010: n2615_o = 1'b0;
      3'b001: n2615_o = 1'b1;
      default: n2615_o = 1'b0;
    endcase
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2618_o = 1'b0;
      3'b010: n2618_o = 1'b1;
      3'b001: n2618_o = 1'b0;
      default: n2618_o = 1'b0;
    endcase
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2620_o = n2595_o;
      3'b010: n2620_o = 1'b0;
      3'b001: n2620_o = 1'b0;
      default: n2620_o = 1'b0;
    endcase
  /* decoder.vhd:905:9  */
  always @*
    case (n2598_o)
      3'b100: n2623_o = 1'b1;
      3'b010: n2623_o = 1'b0;
      3'b001: n2623_o = 1'b0;
      default: n2623_o = 1'b0;
    endcase
  /* decoder.vhd:902:7  */
  assign n2625_o = opc_mnemonic_s == 6'b001100;
  /* decoder.vhd:947:28  */
  assign n2626_o = opc_opcode_q[6];
  /* decoder.vhd:947:13  */
  assign n2629_o = n2626_o ? 1'b1 : 1'b0;
  /* decoder.vhd:947:13  */
  assign n2632_o = n2626_o ? 1'b1 : 1'b0;
  /* decoder.vhd:945:11  */
  assign n2634_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:956:28  */
  assign n2635_o = opc_opcode_q[6];
  /* decoder.vhd:956:32  */
  assign n2636_o = ~n2635_o;
  /* decoder.vhd:956:13  */
  assign n2639_o = n2636_o ? 1'b1 : 1'b0;
  /* decoder.vhd:956:13  */
  assign n2642_o = n2636_o ? 1'b0 : 1'b1;
  /* decoder.vhd:952:11  */
  assign n2644_o = clk_mstate_i == 3'b100;
  assign n2645_o = {n2644_o, n2634_o};
  /* decoder.vhd:944:9  */
  always @*
    case (n2645_o)
      2'b10: n2647_o = n2639_o;
      2'b01: n2647_o = 1'b0;
      default: n2647_o = 1'b0;
    endcase
  /* decoder.vhd:944:9  */
  always @*
    case (n2645_o)
      2'b10: n2649_o = 1'b0;
      2'b01: n2649_o = n2629_o;
      default: n2649_o = 1'b0;
    endcase
  /* decoder.vhd:944:9  */
  always @*
    case (n2645_o)
      2'b10: n2652_o = 1'b1;
      2'b01: n2652_o = 1'b0;
      default: n2652_o = 1'b0;
    endcase
  /* decoder.vhd:944:9  */
  always @*
    case (n2645_o)
      2'b10: n2654_o = 1'b0;
      2'b01: n2654_o = n2632_o;
      default: n2654_o = 1'b0;
    endcase
  /* decoder.vhd:944:9  */
  always @*
    case (n2645_o)
      2'b10: n2657_o = 4'b1000;
      2'b01: n2657_o = 4'b1100;
      default: n2657_o = 4'b1100;
    endcase
  /* decoder.vhd:944:9  */
  always @*
    case (n2645_o)
      2'b10: n2659_o = n2642_o;
      2'b01: n2659_o = 1'b0;
      default: n2659_o = 1'b0;
    endcase
  /* decoder.vhd:943:7  */
  assign n2661_o = opc_mnemonic_s == 6'b001101;
  /* decoder.vhd:971:25  */
  assign n2663_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:972:26  */
  assign n2664_o = opc_opcode_q[4];
  /* decoder.vhd:972:11  */
  assign n2667_o = n2664_o ? 1'b0 : 1'b1;
  /* decoder.vhd:972:11  */
  assign n2670_o = n2664_o ? 1'b1 : 1'b0;
  /* decoder.vhd:971:9  */
  assign n2672_o = n2663_o ? n2667_o : 1'b0;
  /* decoder.vhd:971:9  */
  assign n2674_o = n2663_o ? n2670_o : 1'b0;
  /* decoder.vhd:970:7  */
  assign n2676_o = opc_mnemonic_s == 6'b001110;
  /* decoder.vhd:981:25  */
  assign n2678_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:982:26  */
  assign n2679_o = opc_opcode_q[4];
  /* decoder.vhd:982:11  */
  assign n2682_o = n2679_o ? 1'b0 : 1'b1;
  /* decoder.vhd:982:11  */
  assign n2685_o = n2679_o ? 1'b1 : 1'b0;
  /* decoder.vhd:981:9  */
  assign n2687_o = n2678_o ? n2682_o : 1'b0;
  /* decoder.vhd:981:9  */
  assign n2689_o = n2678_o ? n2685_o : 1'b0;
  /* decoder.vhd:980:7  */
  assign n2691_o = opc_mnemonic_s == 6'b001111;
  /* decoder.vhd:993:12  */
  assign n2692_o = ~clk_second_cycle_i;
  /* decoder.vhd:996:13  */
  assign n2694_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1002:13  */
  assign n2697_o = clk_mstate_i == 3'b100;
  assign n2698_o = {n2697_o, n2694_o};
  /* decoder.vhd:994:11  */
  always @*
    case (n2698_o)
      2'b10: n2701_o = 1'b0;
      2'b01: n2701_o = 1'b1;
      default: n2701_o = 1'b0;
    endcase
  /* decoder.vhd:994:11  */
  always @*
    case (n2698_o)
      2'b10: n2704_o = 1'b1;
      2'b01: n2704_o = 1'b0;
      default: n2704_o = 1'b0;
    endcase
  /* decoder.vhd:994:11  */
  always @*
    case (n2698_o)
      2'b10: n2707_o = 1'b0;
      2'b01: n2707_o = 1'b1;
      default: n2707_o = 1'b0;
    endcase
  /* decoder.vhd:994:11  */
  always @*
    case (n2698_o)
      2'b10: n2710_o = 4'b1000;
      2'b01: n2710_o = 4'b1100;
      default: n2710_o = 4'b1100;
    endcase
  /* decoder.vhd:994:11  */
  always @*
    case (n2698_o)
      2'b10: n2713_o = 1'b1;
      2'b01: n2713_o = 1'b0;
      default: n2713_o = 1'b0;
    endcase
  /* decoder.vhd:994:11  */
  always @*
    case (n2698_o)
      2'b10: n2716_o = 4'b0001;
      2'b01: n2716_o = 4'b0000;
      default: n2716_o = 4'b0000;
    endcase
  assign n2717_o = opc_opcode_q[5];
  /* decoder.vhd:994:11  */
  always @*
    case (n2698_o)
      2'b10: n2718_o = 1'b0;
      2'b01: n2718_o = n2717_o;
      default: n2718_o = n2717_o;
    endcase
  /* decoder.vhd:994:11  */
  always @*
    case (n2698_o)
      2'b10: n2721_o = 1'b1;
      2'b01: n2721_o = 1'b0;
      default: n2721_o = 1'b0;
    endcase
  /* decoder.vhd:1019:27  */
  assign n2723_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1019:37  */
  assign n2724_o = cnd_take_branch_i & n2723_o;
  /* decoder.vhd:1019:11  */
  assign n2730_o = n2724_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1019:11  */
  assign n2733_o = n2724_o ? 1'b1 : 1'b0;
  /* decoder.vhd:993:9  */
  assign n2735_o = n2692_o ? n2701_o : 1'b0;
  /* decoder.vhd:993:9  */
  assign n2737_o = n2692_o ? n2704_o : 1'b0;
  /* decoder.vhd:993:9  */
  assign n2739_o = n2692_o ? n2707_o : 1'b0;
  /* decoder.vhd:993:9  */
  assign n2741_o = n2692_o ? 1'b0 : n2730_o;
  /* decoder.vhd:993:9  */
  assign n2743_o = n2692_o ? n2710_o : 4'b1100;
  /* decoder.vhd:993:9  */
  assign n2745_o = n2692_o ? n2713_o : 1'b0;
  /* decoder.vhd:993:9  */
  assign n2747_o = n2692_o ? n2716_o : 4'b0000;
  assign n2748_o = opc_opcode_q[5];
  /* decoder.vhd:993:9  */
  assign n2749_o = n2692_o ? n2718_o : n2748_o;
  /* decoder.vhd:993:9  */
  assign n2751_o = n2692_o ? 1'b0 : n2733_o;
  /* decoder.vhd:993:9  */
  assign n2753_o = n2692_o ? n2721_o : 1'b0;
  /* decoder.vhd:990:7  */
  assign n2755_o = opc_mnemonic_s == 6'b010000;
  /* decoder.vhd:1027:25  */
  assign n2757_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1027:9  */
  assign n2760_o = n2757_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1026:7  */
  assign n2762_o = opc_mnemonic_s == 6'b010001;
  /* decoder.vhd:1034:48  */
  assign n2764_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1034:31  */
  assign n2765_o = n2764_o & clk_second_cycle_i;
  /* decoder.vhd:1037:26  */
  assign n2766_o = opc_opcode_q[1];
  /* decoder.vhd:1037:30  */
  assign n2767_o = ~n2766_o;
  /* decoder.vhd:1037:11  */
  assign n2770_o = n2767_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1037:11  */
  assign n2773_o = n2767_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1034:9  */
  assign n2776_o = n2765_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1034:9  */
  assign n2778_o = n2765_o ? n2770_o : 1'b0;
  /* decoder.vhd:1034:9  */
  assign n2780_o = n2765_o ? n2773_o : 1'b0;
  /* decoder.vhd:1032:7  */
  assign n2782_o = opc_mnemonic_s == 6'b010010;
  /* decoder.vhd:1049:48  */
  assign n2784_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1049:31  */
  assign n2785_o = n2784_o & clk_second_cycle_i;
  /* decoder.vhd:1049:9  */
  assign n2788_o = n2785_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1049:9  */
  assign n2791_o = n2785_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1045:7  */
  assign n2793_o = opc_mnemonic_s == 6'b010100;
  /* decoder.vhd:1061:28  */
  assign n2794_o = opc_opcode_q[3];
  /* decoder.vhd:1061:32  */
  assign n2795_o = ~n2794_o;
  /* decoder.vhd:1060:44  */
  assign n2797_o = 1'b0 | n2795_o;
  /* decoder.vhd:1060:13  */
  assign n2804_o = n2797_o ? 1'b1 : n2073_o;
  /* decoder.vhd:1060:13  */
  assign n2807_o = n2797_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1060:13  */
  assign n2810_o = n2797_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1059:11  */
  assign n2812_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1067:28  */
  assign n2813_o = opc_opcode_q[3:2];
  /* decoder.vhd:1067:41  */
  assign n2815_o = n2813_o != 2'b01;
  /* decoder.vhd:1067:13  */
  assign n2818_o = n2815_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1067:13  */
  assign n2821_o = n2815_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1065:11  */
  assign n2823_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1076:28  */
  assign n2824_o = opc_opcode_q[3:2];
  /* decoder.vhd:1076:41  */
  assign n2826_o = n2824_o == 2'b01;
  /* decoder.vhd:1076:13  */
  assign n2829_o = n2826_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1076:13  */
  assign n2832_o = n2826_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1072:11  */
  assign n2834_o = clk_mstate_i == 3'b100;
  assign n2835_o = {n2834_o, n2823_o, n2812_o};
  /* decoder.vhd:1057:9  */
  always @*
    case (n2835_o)
      3'b100: n2837_o = n2829_o;
      3'b010: n2837_o = 1'b0;
      3'b001: n2837_o = 1'b0;
      default: n2837_o = 1'b0;
    endcase
  /* decoder.vhd:1057:9  */
  always @*
    case (n2835_o)
      3'b100: n2839_o = 1'b0;
      3'b010: n2839_o = n2818_o;
      3'b001: n2839_o = 1'b0;
      default: n2839_o = 1'b0;
    endcase
  /* decoder.vhd:1057:9  */
  always @*
    case (n2835_o)
      3'b100: n2842_o = 1'b1;
      3'b010: n2842_o = 1'b0;
      3'b001: n2842_o = 1'b0;
      default: n2842_o = 1'b0;
    endcase
  /* decoder.vhd:1057:9  */
  always @*
    case (n2835_o)
      3'b100: n2843_o = n2073_o;
      3'b010: n2843_o = n2073_o;
      3'b001: n2843_o = n2804_o;
      default: n2843_o = n2073_o;
    endcase
  /* decoder.vhd:1057:9  */
  always @*
    case (n2835_o)
      3'b100: n2845_o = 1'b0;
      3'b010: n2845_o = n2821_o;
      3'b001: n2845_o = n2807_o;
      default: n2845_o = 1'b0;
    endcase
  /* decoder.vhd:1057:9  */
  always @*
    case (n2835_o)
      3'b100: n2848_o = 4'b1001;
      3'b010: n2848_o = 4'b1100;
      3'b001: n2848_o = 4'b1100;
      default: n2848_o = 4'b1100;
    endcase
  /* decoder.vhd:1057:9  */
  always @*
    case (n2835_o)
      3'b100: n2850_o = 2'b01;
      3'b010: n2850_o = 2'b01;
      3'b001: n2850_o = n2810_o;
      default: n2850_o = 2'b01;
    endcase
  /* decoder.vhd:1057:9  */
  always @*
    case (n2835_o)
      3'b100: n2852_o = n2832_o;
      3'b010: n2852_o = 1'b0;
      3'b001: n2852_o = 1'b0;
      default: n2852_o = 1'b0;
    endcase
  /* decoder.vhd:1056:7  */
  assign n2854_o = opc_mnemonic_s == 6'b010011;
  /* decoder.vhd:1094:12  */
  assign n2855_o = ~clk_second_cycle_i;
  /* decoder.vhd:1096:27  */
  assign n2857_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1096:11  */
  assign n2860_o = n2857_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1096:11  */
  assign n2863_o = n2857_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1105:27  */
  assign n2865_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1105:37  */
  assign n2866_o = cnd_take_branch_i & n2865_o;
  /* decoder.vhd:1105:11  */
  assign n2872_o = n2866_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1105:11  */
  assign n2875_o = n2866_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1094:9  */
  assign n2877_o = n2855_o ? n2860_o : 1'b0;
  /* decoder.vhd:1094:9  */
  assign n2879_o = n2855_o ? 1'b0 : n2872_o;
  /* decoder.vhd:1094:9  */
  assign n2881_o = n2855_o ? n2863_o : 1'b0;
  /* decoder.vhd:1094:9  */
  assign n2883_o = n2855_o ? 1'b0 : n2875_o;
  /* decoder.vhd:1090:7  */
  assign n2885_o = opc_mnemonic_s == 6'b010101;
  /* decoder.vhd:1116:12  */
  assign n2886_o = ~clk_second_cycle_i;
  /* decoder.vhd:1118:27  */
  assign n2888_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1120:48  */
  assign n2889_o = opc_opcode_q[4];
  /* decoder.vhd:1118:11  */
  assign n2892_o = n2888_o ? 1'b1 : 1'b0;
  assign n2893_o = opc_opcode_q[5];
  /* decoder.vhd:1116:9  */
  assign n2894_o = n2912_o ? n2889_o : n2893_o;
  /* decoder.vhd:1126:27  */
  assign n2896_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1126:37  */
  assign n2897_o = cnd_take_branch_i & n2896_o;
  /* decoder.vhd:1126:11  */
  assign n2903_o = n2897_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1126:11  */
  assign n2906_o = n2897_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1116:9  */
  assign n2908_o = n2886_o ? 1'b0 : n2903_o;
  /* decoder.vhd:1116:9  */
  assign n2910_o = n2886_o ? n2892_o : 1'b0;
  /* decoder.vhd:1116:9  */
  assign n2912_o = n2886_o & n2888_o;
  /* decoder.vhd:1116:9  */
  assign n2914_o = n2886_o ? 1'b0 : n2906_o;
  /* decoder.vhd:1112:7  */
  assign n2916_o = opc_mnemonic_s == 6'b010110;
  /* decoder.vhd:1136:12  */
  assign n2917_o = ~clk_second_cycle_i;
  /* decoder.vhd:1138:27  */
  assign n2919_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1140:28  */
  assign n2920_o = opc_opcode_q[7];
  /* decoder.vhd:1140:13  */
  assign n2923_o = n2920_o ? 4'b0011 : 4'b0100;
  /* decoder.vhd:1138:11  */
  assign n2926_o = n2919_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1138:11  */
  assign n2928_o = n2919_o ? n2923_o : 4'b0000;
  /* decoder.vhd:1153:27  */
  assign n2930_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1153:37  */
  assign n2931_o = cnd_take_branch_i & n2930_o;
  /* decoder.vhd:1153:11  */
  assign n2937_o = n2931_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1153:11  */
  assign n2940_o = n2931_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1136:9  */
  assign n2942_o = n2917_o ? 1'b0 : n2937_o;
  /* decoder.vhd:1136:9  */
  assign n2944_o = n2917_o ? n2926_o : 1'b0;
  /* decoder.vhd:1136:9  */
  assign n2946_o = n2917_o ? n2928_o : 4'b0000;
  /* decoder.vhd:1136:9  */
  assign n2948_o = n2917_o ? 1'b0 : n2940_o;
  /* decoder.vhd:1133:7  */
  assign n2950_o = opc_mnemonic_s == 6'b010111;
  /* decoder.vhd:1167:13  */
  assign n2952_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1173:40  */
  assign n2954_o = {4'b0000, n2058_o};
  /* decoder.vhd:1173:61  */
  assign n2955_o = opc_opcode_q[7:5];
  /* decoder.vhd:1173:47  */
  assign n2956_o = {n2954_o, n2955_o};
  /* decoder.vhd:1172:13  */
  assign n2958_o = clk_mstate_i == 3'b001;
  assign n2959_o = {n2958_o, n2952_o};
  /* decoder.vhd:1165:11  */
  always @*
    case (n2959_o)
      2'b10: n2962_o = 1'b0;
      2'b01: n2962_o = 1'b1;
      default: n2962_o = 1'b0;
    endcase
  /* decoder.vhd:1165:11  */
  always @*
    case (n2959_o)
      2'b10: n2965_o = 1'b1;
      2'b01: n2965_o = 1'b0;
      default: n2965_o = 1'b0;
    endcase
  /* decoder.vhd:1165:11  */
  always @*
    case (n2959_o)
      2'b10: n2968_o = 1'b0;
      2'b01: n2968_o = 1'b1;
      default: n2968_o = 1'b0;
    endcase
  /* decoder.vhd:1165:11  */
  always @*
    case (n2959_o)
      2'b10: n2969_o = n2956_o;
      2'b01: n2969_o = n2077_o;
      default: n2969_o = n2077_o;
    endcase
  /* decoder.vhd:1165:11  */
  always @*
    case (n2959_o)
      2'b10: n2971_o = 1'b1;
      2'b01: n2971_o = n2081_o;
      default: n2971_o = n2081_o;
    endcase
  /* decoder.vhd:1164:9  */
  assign n2973_o = clk_second_cycle_i ? n2962_o : 1'b0;
  /* decoder.vhd:1164:9  */
  assign n2975_o = clk_second_cycle_i ? n2965_o : 1'b0;
  /* decoder.vhd:1164:9  */
  assign n2977_o = clk_second_cycle_i ? n2968_o : 1'b0;
  /* decoder.vhd:1164:9  */
  assign n2978_o = clk_second_cycle_i ? n2969_o : n2077_o;
  /* decoder.vhd:1164:9  */
  assign n2979_o = clk_second_cycle_i ? n2971_o : n2081_o;
  /* decoder.vhd:1161:7  */
  assign n2981_o = opc_mnemonic_s == 6'b011000;
  /* decoder.vhd:1188:12  */
  assign n2982_o = ~clk_second_cycle_i;
  /* decoder.vhd:1191:27  */
  assign n2984_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1191:11  */
  assign n2987_o = n2984_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1191:11  */
  assign n2990_o = n2984_o ? 2'b01 : 2'b00;
  /* decoder.vhd:1197:27  */
  assign n2992_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1197:11  */
  assign n2995_o = n2992_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1197:11  */
  assign n2998_o = n2992_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1188:9  */
  assign n3000_o = n2982_o ? n2987_o : 1'b0;
  /* decoder.vhd:1188:9  */
  assign n3002_o = n2982_o ? 1'b0 : n2995_o;
  /* decoder.vhd:1188:9  */
  assign n3004_o = n2982_o ? n2990_o : 2'b00;
  /* decoder.vhd:1188:9  */
  assign n3006_o = n2982_o ? 1'b0 : n2998_o;
  /* decoder.vhd:1185:7  */
  assign n3008_o = opc_mnemonic_s == 6'b011001;
  /* decoder.vhd:1210:12  */
  assign n3009_o = ~clk_second_cycle_i;
  /* decoder.vhd:1212:27  */
  assign n3011_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1212:11  */
  assign n3014_o = n3011_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1219:27  */
  assign n3016_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1219:37  */
  assign n3017_o = cnd_take_branch_i & n3016_o;
  /* decoder.vhd:1219:11  */
  assign n3023_o = n3017_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1219:11  */
  assign n3026_o = n3017_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1210:9  */
  assign n3028_o = n3009_o ? 1'b0 : n3023_o;
  /* decoder.vhd:1210:9  */
  assign n3030_o = n3009_o ? n3014_o : 1'b0;
  /* decoder.vhd:1210:9  */
  assign n3032_o = n3009_o ? 1'b0 : n3026_o;
  /* decoder.vhd:1206:7  */
  assign n3034_o = opc_mnemonic_s == 6'b011010;
  /* decoder.vhd:1228:24  */
  assign n3035_o = opc_opcode_q[6];
  /* decoder.vhd:1228:28  */
  assign n3036_o = ~n3035_o;
  /* decoder.vhd:1228:9  */
  assign n3039_o = n3036_o ? 4'b0110 : 4'b0111;
  /* decoder.vhd:1234:12  */
  assign n3040_o = ~clk_second_cycle_i;
  /* decoder.vhd:1236:27  */
  assign n3042_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1238:48  */
  assign n3043_o = opc_opcode_q[4];
  /* decoder.vhd:1236:11  */
  assign n3046_o = n3042_o ? 1'b1 : 1'b0;
  assign n3047_o = opc_opcode_q[5];
  /* decoder.vhd:1234:9  */
  assign n3048_o = n3066_o ? n3043_o : n3047_o;
  /* decoder.vhd:1244:27  */
  assign n3050_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1244:37  */
  assign n3051_o = cnd_take_branch_i & n3050_o;
  /* decoder.vhd:1244:11  */
  assign n3057_o = n3051_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1244:11  */
  assign n3060_o = n3051_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1234:9  */
  assign n3062_o = n3040_o ? 1'b0 : n3057_o;
  /* decoder.vhd:1234:9  */
  assign n3064_o = n3040_o ? n3046_o : 1'b0;
  /* decoder.vhd:1234:9  */
  assign n3066_o = n3040_o & n3042_o;
  /* decoder.vhd:1234:9  */
  assign n3068_o = n3040_o ? 1'b0 : n3060_o;
  /* decoder.vhd:1226:7  */
  assign n3070_o = opc_mnemonic_s == 6'b011011;
  /* decoder.vhd:1255:12  */
  assign n3071_o = ~clk_second_cycle_i;
  /* decoder.vhd:1257:27  */
  assign n3073_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1257:11  */
  assign n3076_o = n3073_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1257:11  */
  assign n3079_o = n3073_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1265:27  */
  assign n3081_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1265:37  */
  assign n3082_o = cnd_take_branch_i & n3081_o;
  /* decoder.vhd:1265:11  */
  assign n3088_o = n3082_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1265:11  */
  assign n3091_o = n3082_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1255:9  */
  assign n3093_o = n3071_o ? 1'b0 : n3088_o;
  /* decoder.vhd:1255:9  */
  assign n3095_o = n3071_o ? n3076_o : 1'b0;
  /* decoder.vhd:1255:9  */
  assign n3097_o = n3071_o ? 1'b0 : n3091_o;
  /* decoder.vhd:1255:9  */
  assign n3099_o = n3071_o ? n3079_o : 1'b0;
  /* decoder.vhd:1251:7  */
  assign n3101_o = opc_mnemonic_s == 6'b011100;
  /* decoder.vhd:1276:12  */
  assign n3102_o = ~clk_second_cycle_i;
  /* decoder.vhd:1278:27  */
  assign n3104_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1281:48  */
  assign n3105_o = opc_opcode_q[6];
  /* decoder.vhd:1278:11  */
  assign n3108_o = n3104_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1278:11  */
  assign n3111_o = n3104_o ? 1'b1 : 1'b0;
  assign n3112_o = opc_opcode_q[5];
  /* decoder.vhd:1276:9  */
  assign n3113_o = n3133_o ? n3105_o : n3112_o;
  /* decoder.vhd:1287:27  */
  assign n3115_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1287:37  */
  assign n3116_o = cnd_take_branch_i & n3115_o;
  /* decoder.vhd:1287:11  */
  assign n3122_o = n3116_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1287:11  */
  assign n3125_o = n3116_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1276:9  */
  assign n3127_o = n3102_o ? n3108_o : 1'b0;
  /* decoder.vhd:1276:9  */
  assign n3129_o = n3102_o ? 1'b0 : n3122_o;
  /* decoder.vhd:1276:9  */
  assign n3131_o = n3102_o ? n3111_o : 1'b0;
  /* decoder.vhd:1276:9  */
  assign n3133_o = n3102_o & n3104_o;
  /* decoder.vhd:1276:9  */
  assign n3135_o = n3102_o ? 1'b0 : n3125_o;
  /* decoder.vhd:1272:7  */
  assign n3137_o = opc_mnemonic_s == 6'b011101;
  /* decoder.vhd:1299:48  */
  assign n3139_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1299:31  */
  assign n3140_o = n3139_o & clk_second_cycle_i;
  /* decoder.vhd:1299:9  */
  assign n3143_o = n3140_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1294:7  */
  assign n3145_o = opc_mnemonic_s == 6'b011110;
  /* decoder.vhd:1309:28  */
  assign n3146_o = opc_opcode_q[3];
  /* decoder.vhd:1309:32  */
  assign n3147_o = ~n3146_o;
  /* decoder.vhd:1308:44  */
  assign n3149_o = 1'b0 | n3147_o;
  /* decoder.vhd:1308:13  */
  assign n3156_o = n3149_o ? 1'b1 : n2073_o;
  /* decoder.vhd:1308:13  */
  assign n3159_o = n3149_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1308:13  */
  assign n3162_o = n3149_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1307:11  */
  assign n3164_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1314:11  */
  assign n3169_o = clk_mstate_i == 3'b011;
  assign n3170_o = {n3169_o, n3164_o};
  /* decoder.vhd:1305:9  */
  always @*
    case (n3170_o)
      2'b10: n3173_o = 1'b1;
      2'b01: n3173_o = 1'b0;
      default: n3173_o = 1'b0;
    endcase
  /* decoder.vhd:1305:9  */
  always @*
    case (n3170_o)
      2'b10: n3176_o = 1'b1;
      2'b01: n3176_o = 1'b0;
      default: n3176_o = 1'b0;
    endcase
  /* decoder.vhd:1305:9  */
  always @*
    case (n3170_o)
      2'b10: n3177_o = n2073_o;
      2'b01: n3177_o = n3156_o;
      default: n3177_o = n2073_o;
    endcase
  /* decoder.vhd:1305:9  */
  always @*
    case (n3170_o)
      2'b10: n3180_o = 1'b1;
      2'b01: n3180_o = n3159_o;
      default: n3180_o = 1'b0;
    endcase
  /* decoder.vhd:1305:9  */
  always @*
    case (n3170_o)
      2'b10: n3182_o = 2'b01;
      2'b01: n3182_o = n3162_o;
      default: n3182_o = 2'b01;
    endcase
  /* decoder.vhd:1304:7  */
  assign n3184_o = opc_mnemonic_s == 6'b100000;
  /* decoder.vhd:1325:25  */
  assign n3186_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1325:9  */
  assign n3189_o = n3186_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1325:9  */
  assign n3192_o = n3186_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1325:9  */
  assign n3195_o = n3186_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1324:7  */
  assign n3197_o = opc_mnemonic_s == 6'b011111;
  /* decoder.vhd:1333:25  */
  assign n3199_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1333:9  */
  assign n3202_o = n3199_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1333:9  */
  assign n3205_o = n3199_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1333:9  */
  assign n3208_o = n3199_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1332:7  */
  assign n3210_o = opc_mnemonic_s == 6'b100001;
  /* decoder.vhd:1345:28  */
  assign n3211_o = opc_opcode_q[3];
  /* decoder.vhd:1345:32  */
  assign n3212_o = ~n3211_o;
  /* decoder.vhd:1344:44  */
  assign n3214_o = 1'b0 | n3212_o;
  /* decoder.vhd:1344:13  */
  assign n3221_o = n3214_o ? 1'b1 : n2073_o;
  /* decoder.vhd:1344:13  */
  assign n3224_o = n3214_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1344:13  */
  assign n3227_o = n3214_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1343:11  */
  assign n3229_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1350:11  */
  assign n3231_o = clk_mstate_i == 3'b100;
  assign n3232_o = {n3231_o, n3229_o};
  /* decoder.vhd:1341:9  */
  always @*
    case (n3232_o)
      2'b10: n3235_o = 1'b1;
      2'b01: n3235_o = 1'b0;
      default: n3235_o = 1'b0;
    endcase
  /* decoder.vhd:1341:9  */
  always @*
    case (n3232_o)
      2'b10: n3236_o = n2073_o;
      2'b01: n3236_o = n3221_o;
      default: n3236_o = n2073_o;
    endcase
  /* decoder.vhd:1341:9  */
  always @*
    case (n3232_o)
      2'b10: n3238_o = 1'b0;
      2'b01: n3238_o = n3224_o;
      default: n3238_o = 1'b0;
    endcase
  /* decoder.vhd:1341:9  */
  always @*
    case (n3232_o)
      2'b10: n3240_o = 2'b01;
      2'b01: n3240_o = n3227_o;
      default: n3240_o = 2'b01;
    endcase
  /* decoder.vhd:1341:9  */
  always @*
    case (n3232_o)
      2'b10: n3243_o = 1'b1;
      2'b01: n3243_o = 1'b0;
      default: n3243_o = 1'b0;
    endcase
  /* decoder.vhd:1340:7  */
  assign n3245_o = opc_mnemonic_s == 6'b100010;
  /* decoder.vhd:1364:12  */
  assign n3246_o = ~clk_second_cycle_i;
  /* decoder.vhd:1364:52  */
  assign n3248_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1364:35  */
  assign n3249_o = n3248_o & n3246_o;
  /* decoder.vhd:1366:26  */
  assign n3250_o = opc_opcode_q[3];
  /* decoder.vhd:1366:30  */
  assign n3251_o = ~n3250_o;
  /* decoder.vhd:1365:42  */
  assign n3253_o = 1'b0 | n3251_o;
  /* decoder.vhd:1364:9  */
  assign n3260_o = n3267_o ? 1'b1 : n2073_o;
  /* decoder.vhd:1365:11  */
  assign n3263_o = n3253_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1365:11  */
  assign n3266_o = n3253_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1364:9  */
  assign n3267_o = n3249_o & n3253_o;
  /* decoder.vhd:1364:9  */
  assign n3269_o = n3249_o ? n3263_o : 1'b0;
  /* decoder.vhd:1364:9  */
  assign n3271_o = n3249_o ? n3266_o : 2'b01;
  /* decoder.vhd:1373:48  */
  assign n3273_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1373:31  */
  assign n3274_o = n3273_o & clk_second_cycle_i;
  /* decoder.vhd:1373:9  */
  assign n3277_o = n3274_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1360:7  */
  assign n3279_o = opc_mnemonic_s == 6'b100011;
  /* decoder.vhd:1379:25  */
  assign n3281_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1380:26  */
  assign n3282_o = opc_opcode_q[5];
  /* decoder.vhd:1380:11  */
  assign n3285_o = n3282_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1380:11  */
  assign n3288_o = n3282_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1380:11  */
  assign n3291_o = n3282_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1380:11  */
  assign n3294_o = n3282_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1379:9  */
  assign n3296_o = n3281_o ? n3285_o : 1'b0;
  /* decoder.vhd:1379:9  */
  assign n3298_o = n3281_o ? n3288_o : 1'b0;
  /* decoder.vhd:1379:9  */
  assign n3300_o = n3281_o ? n3291_o : 1'b0;
  /* decoder.vhd:1379:9  */
  assign n3302_o = n3281_o ? n3294_o : 1'b0;
  /* decoder.vhd:1378:7  */
  assign n3304_o = opc_mnemonic_s == 6'b100100;
  /* decoder.vhd:1393:12  */
  assign n3305_o = ~clk_second_cycle_i;
  /* decoder.vhd:1399:53  */
  assign n3307_o = opc_opcode_q[1:0];
  /* decoder.vhd:1401:32  */
  assign n3308_o = opc_opcode_q[7:4];
  /* decoder.vhd:1402:17  */
  assign n3311_o = n3308_o == 4'b1001;
  /* decoder.vhd:1404:17  */
  assign n3314_o = n3308_o == 4'b1000;
  /* decoder.vhd:1406:17  */
  assign n3317_o = n3308_o == 4'b0011;
  assign n3318_o = {n3317_o, n3314_o, n3311_o};
  assign n3319_o = n2075_o[3:2];
  assign n3320_o = n2076_o[3:2];
  /* decoder.vhd:593:5  */
  assign n3321_o = n2062_o ? n3319_o : n3320_o;
  /* decoder.vhd:1401:15  */
  always @*
    case (n3318_o)
      3'b100: n3322_o = 2'b01;
      3'b010: n3322_o = 2'b10;
      3'b001: n3322_o = 2'b11;
      default: n3322_o = n3321_o;
    endcase
  /* decoder.vhd:1396:13  */
  assign n3324_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1417:13  */
  assign n3326_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1423:13  */
  assign n3328_o = clk_mstate_i == 3'b100;
  assign n3329_o = {n3328_o, n3326_o, n3324_o};
  /* decoder.vhd:1394:11  */
  always @*
    case (n3329_o)
      3'b100: n3332_o = 1'b0;
      3'b010: n3332_o = 1'b1;
      3'b001: n3332_o = 1'b0;
      default: n3332_o = 1'b0;
    endcase
  /* decoder.vhd:1394:11  */
  always @*
    case (n3329_o)
      3'b100: n3336_o = 1'b0;
      3'b010: n3336_o = 1'b1;
      3'b001: n3336_o = 1'b1;
      default: n3336_o = 1'b0;
    endcase
  assign n3337_o = n2075_o[1:0];
  assign n3338_o = n2076_o[1:0];
  /* decoder.vhd:593:5  */
  assign n3339_o = n2062_o ? n3337_o : n3338_o;
  /* decoder.vhd:1394:11  */
  always @*
    case (n3329_o)
      3'b100: n3340_o = n3339_o;
      3'b010: n3340_o = n3339_o;
      3'b001: n3340_o = n3307_o;
      default: n3340_o = n3339_o;
    endcase
  assign n3341_o = n2075_o[3:2];
  assign n3342_o = n2076_o[3:2];
  /* decoder.vhd:593:5  */
  assign n3343_o = n2062_o ? n3341_o : n3342_o;
  /* decoder.vhd:1394:11  */
  always @*
    case (n3329_o)
      3'b100: n3344_o = n3343_o;
      3'b010: n3344_o = n3343_o;
      3'b001: n3344_o = n3322_o;
      default: n3344_o = n3343_o;
    endcase
  assign n3345_o = n2075_o[7:4];
  assign n3346_o = n2076_o[7:4];
  /* decoder.vhd:593:5  */
  assign n3347_o = n2062_o ? n3345_o : n3346_o;
  /* decoder.vhd:1394:11  */
  always @*
    case (n3329_o)
      3'b100: n3348_o = n3347_o;
      3'b010: n3348_o = n3347_o;
      3'b001: n3348_o = 4'b0000;
      default: n3348_o = n3347_o;
    endcase
  /* decoder.vhd:1394:11  */
  always @*
    case (n3329_o)
      3'b100: n3350_o = n2081_o;
      3'b010: n3350_o = n2081_o;
      3'b001: n3350_o = 1'b1;
      default: n3350_o = n2081_o;
    endcase
  /* decoder.vhd:1394:11  */
  always @*
    case (n3329_o)
      3'b100: n3354_o = 1'b1;
      3'b010: n3354_o = 1'b1;
      3'b001: n3354_o = 1'b0;
      default: n3354_o = 1'b0;
    endcase
  /* decoder.vhd:1433:27  */
  assign n3356_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1433:53  */
  assign n3358_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1433:37  */
  assign n3359_o = n3356_o | n3358_o;
  /* decoder.vhd:1433:11  */
  assign n3362_o = n3359_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1393:9  */
  assign n3364_o = n3305_o ? n3332_o : 1'b0;
  /* decoder.vhd:1393:9  */
  assign n3366_o = n3305_o ? n3336_o : 1'b0;
  assign n3367_o = {n3348_o, n3344_o, n3340_o};
  /* decoder.vhd:1393:9  */
  assign n3368_o = n3305_o ? n3367_o : n2077_o;
  /* decoder.vhd:1393:9  */
  assign n3369_o = n3305_o ? n3350_o : n2081_o;
  /* decoder.vhd:1393:9  */
  assign n3370_o = n3305_o ? n3354_o : n3362_o;
  /* decoder.vhd:1390:7  */
  assign n3372_o = opc_mnemonic_s == 6'b101100;
  /* decoder.vhd:1443:12  */
  assign n3373_o = ~clk_second_cycle_i;
  /* decoder.vhd:1449:53  */
  assign n3374_o = opc_opcode_q[1:0];
  /* decoder.vhd:1448:48  */
  assign n3376_o = {6'b000000, n3374_o};
  /* decoder.vhd:1446:13  */
  assign n3378_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1455:13  */
  assign n3381_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1462:13  */
  assign n3383_o = clk_mstate_i == 3'b100;
  assign n3384_o = {n3383_o, n3381_o, n3378_o};
  /* decoder.vhd:1444:11  */
  always @*
    case (n3384_o)
      3'b100: n3388_o = 1'b0;
      3'b010: n3388_o = 1'b1;
      3'b001: n3388_o = 1'b1;
      default: n3388_o = 1'b0;
    endcase
  assign n3389_o = n3376_o[3:0];
  assign n3390_o = n2075_o[3:0];
  assign n3391_o = n2076_o[3:0];
  /* decoder.vhd:593:5  */
  assign n3392_o = n2062_o ? n3390_o : n3391_o;
  /* decoder.vhd:1444:11  */
  always @*
    case (n3384_o)
      3'b100: n3393_o = n3392_o;
      3'b010: n3393_o = 4'b1111;
      3'b001: n3393_o = n3389_o;
      default: n3393_o = n3392_o;
    endcase
  assign n3394_o = n3376_o[7:4];
  assign n3395_o = n2075_o[7:4];
  assign n3396_o = n2076_o[7:4];
  /* decoder.vhd:593:5  */
  assign n3397_o = n2062_o ? n3395_o : n3396_o;
  /* decoder.vhd:1444:11  */
  always @*
    case (n3384_o)
      3'b100: n3398_o = n3397_o;
      3'b010: n3398_o = n3397_o;
      3'b001: n3398_o = n3394_o;
      default: n3398_o = n3397_o;
    endcase
  /* decoder.vhd:1444:11  */
  always @*
    case (n3384_o)
      3'b100: n3401_o = n2081_o;
      3'b010: n3401_o = 1'b1;
      3'b001: n3401_o = 1'b1;
      default: n3401_o = n2081_o;
    endcase
  /* decoder.vhd:1444:11  */
  always @*
    case (n3384_o)
      3'b100: n3405_o = 1'b1;
      3'b010: n3405_o = 1'b1;
      3'b001: n3405_o = 1'b0;
      default: n3405_o = 1'b0;
    endcase
  /* decoder.vhd:1473:13  */
  assign n3407_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1478:13  */
  assign n3409_o = clk_mstate_i == 3'b001;
  assign n3410_o = {n3409_o, n3407_o};
  /* decoder.vhd:1471:11  */
  always @*
    case (n3410_o)
      2'b10: n3413_o = 1'b1;
      2'b01: n3413_o = 1'b0;
      default: n3413_o = 1'b0;
    endcase
  /* decoder.vhd:1471:11  */
  always @*
    case (n3410_o)
      2'b10: n3416_o = 1'b1;
      2'b01: n3416_o = 1'b0;
      default: n3416_o = 1'b0;
    endcase
  /* decoder.vhd:1471:11  */
  always @*
    case (n3410_o)
      2'b10: n3419_o = 1'b1;
      2'b01: n3419_o = 1'b0;
      default: n3419_o = 1'b0;
    endcase
  /* decoder.vhd:1471:11  */
  always @*
    case (n3410_o)
      2'b10: n3423_o = 1'b1;
      2'b01: n3423_o = 1'b1;
      default: n3423_o = 1'b0;
    endcase
  /* decoder.vhd:1443:9  */
  assign n3425_o = n3373_o ? 1'b0 : n3413_o;
  /* decoder.vhd:1443:9  */
  assign n3427_o = n3373_o ? n3388_o : 1'b0;
  /* decoder.vhd:1443:9  */
  assign n3429_o = n3373_o ? 1'b0 : n3416_o;
  /* decoder.vhd:1443:9  */
  assign n3431_o = n3373_o ? 1'b0 : n3419_o;
  assign n3432_o = {n3398_o, n3393_o};
  /* decoder.vhd:1443:9  */
  assign n3433_o = n3373_o ? n3432_o : n2077_o;
  /* decoder.vhd:1443:9  */
  assign n3434_o = n3373_o ? n3401_o : n2081_o;
  /* decoder.vhd:1443:9  */
  assign n3435_o = n3373_o ? n3405_o : n3423_o;
  /* decoder.vhd:1440:7  */
  assign n3437_o = opc_mnemonic_s == 6'b100101;
  /* decoder.vhd:1495:12  */
  assign n3438_o = ~clk_second_cycle_i;
  /* decoder.vhd:1498:27  */
  assign n3440_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1500:28  */
  assign n3441_o = opc_opcode_q[6];
  /* decoder.vhd:1500:32  */
  assign n3442_o = ~n3441_o;
  /* decoder.vhd:1500:13  */
  assign n3445_o = n3442_o ? 2'b01 : 2'b10;
  /* decoder.vhd:1498:11  */
  assign n3448_o = n3440_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1498:11  */
  assign n3450_o = n3440_o ? n3445_o : 2'b00;
  /* decoder.vhd:1508:27  */
  assign n3452_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1508:11  */
  assign n3455_o = n3452_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1508:11  */
  assign n3458_o = n3452_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1495:9  */
  assign n3460_o = n3438_o ? 1'b0 : n3455_o;
  /* decoder.vhd:1495:9  */
  assign n3462_o = n3438_o ? n3448_o : 1'b0;
  /* decoder.vhd:1495:9  */
  assign n3464_o = n3438_o ? n3450_o : 2'b00;
  /* decoder.vhd:1495:9  */
  assign n3466_o = n3438_o ? 1'b0 : n3458_o;
  /* decoder.vhd:1492:7  */
  assign n3468_o = opc_mnemonic_s == 6'b100110;
  /* decoder.vhd:1522:24  */
  assign n3469_o = opc_opcode_q[4];
  /* decoder.vhd:1522:28  */
  assign n3470_o = ~n3469_o;
  /* decoder.vhd:1522:9  */
  assign n3473_o = n3470_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1522:9  */
  assign n3476_o = n3470_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1528:12  */
  assign n3477_o = ~clk_second_cycle_i;
  /* decoder.vhd:1532:13  */
  assign n3479_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1538:30  */
  assign n3480_o = opc_opcode_q[4];
  /* decoder.vhd:1538:15  */
  assign n3483_o = n3480_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1538:15  */
  assign n3486_o = n3480_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1537:13  */
  assign n3488_o = clk_mstate_i == 3'b100;
  assign n3489_o = {n3488_o, n3479_o};
  /* decoder.vhd:1530:11  */
  always @*
    case (n3489_o)
      2'b10: n3491_o = n3483_o;
      2'b01: n3491_o = 1'b0;
      default: n3491_o = 1'b0;
    endcase
  /* decoder.vhd:1530:11  */
  always @*
    case (n3489_o)
      2'b10: n3494_o = n3486_o;
      2'b01: n3494_o = 1'b1;
      default: n3494_o = 1'b0;
    endcase
  /* decoder.vhd:1530:11  */
  always @*
    case (n3489_o)
      2'b10: n3497_o = 1'b0;
      2'b01: n3497_o = 1'b1;
      default: n3497_o = 1'b0;
    endcase
  /* decoder.vhd:1548:27  */
  assign n3499_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1549:28  */
  assign n3500_o = opc_opcode_q[4];
  /* decoder.vhd:1549:32  */
  assign n3501_o = ~n3500_o;
  /* decoder.vhd:1549:13  */
  assign n3504_o = n3501_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1549:13  */
  assign n3507_o = n3501_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1549:13  */
  assign n3510_o = n3501_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1549:13  */
  assign n3513_o = n3501_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1548:11  */
  assign n3515_o = n3499_o ? n3504_o : 1'b0;
  /* decoder.vhd:1548:11  */
  assign n3517_o = n3499_o ? n3507_o : 1'b0;
  /* decoder.vhd:1548:11  */
  assign n3519_o = n3499_o ? n3510_o : 1'b0;
  /* decoder.vhd:1548:11  */
  assign n3521_o = n3499_o ? n3513_o : 1'b0;
  /* decoder.vhd:1528:9  */
  assign n3523_o = n3477_o ? 1'b0 : n3515_o;
  /* decoder.vhd:1528:9  */
  assign n3524_o = n3477_o ? n3491_o : n3517_o;
  /* decoder.vhd:1528:9  */
  assign n3525_o = n3477_o ? n3494_o : n3519_o;
  /* decoder.vhd:1528:9  */
  assign n3527_o = n3477_o ? n3497_o : 1'b0;
  /* decoder.vhd:1528:9  */
  assign n3529_o = n3477_o ? 1'b0 : n3521_o;
  /* decoder.vhd:1528:9  */
  assign n3532_o = n3477_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1519:7  */
  assign n3534_o = opc_mnemonic_s == 6'b100111;
  /* decoder.vhd:1564:7  */
  assign n3536_o = opc_mnemonic_s == 6'b101000;
  /* decoder.vhd:1573:28  */
  assign n3537_o = opc_opcode_q[3];
  /* decoder.vhd:1573:32  */
  assign n3538_o = ~n3537_o;
  /* decoder.vhd:1572:44  */
  assign n3540_o = 1'b0 | n3538_o;
  /* decoder.vhd:1572:13  */
  assign n3547_o = n3540_o ? 1'b1 : n2073_o;
  /* decoder.vhd:1572:13  */
  assign n3550_o = n3540_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1572:13  */
  assign n3553_o = n3540_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1571:11  */
  assign n3555_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1578:11  */
  assign n3560_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1582:11  */
  assign n3565_o = clk_mstate_i == 3'b100;
  assign n3566_o = {n3565_o, n3560_o, n3555_o};
  /* decoder.vhd:1569:9  */
  always @*
    case (n3566_o)
      3'b100: n3569_o = 1'b1;
      3'b010: n3569_o = 1'b0;
      3'b001: n3569_o = 1'b0;
      default: n3569_o = 1'b0;
    endcase
  /* decoder.vhd:1569:9  */
  always @*
    case (n3566_o)
      3'b100: n3572_o = 1'b0;
      3'b010: n3572_o = 1'b1;
      3'b001: n3572_o = 1'b0;
      default: n3572_o = 1'b0;
    endcase
  /* decoder.vhd:1569:9  */
  always @*
    case (n3566_o)
      3'b100: n3575_o = 1'b1;
      3'b010: n3575_o = 1'b0;
      3'b001: n3575_o = 1'b0;
      default: n3575_o = 1'b0;
    endcase
  /* decoder.vhd:1569:9  */
  always @*
    case (n3566_o)
      3'b100: n3576_o = n2073_o;
      3'b010: n3576_o = n2073_o;
      3'b001: n3576_o = n3547_o;
      default: n3576_o = n2073_o;
    endcase
  /* decoder.vhd:1569:9  */
  always @*
    case (n3566_o)
      3'b100: n3579_o = 1'b0;
      3'b010: n3579_o = 1'b1;
      3'b001: n3579_o = n3550_o;
      default: n3579_o = 1'b0;
    endcase
  /* decoder.vhd:1569:9  */
  always @*
    case (n3566_o)
      3'b100: n3582_o = 4'b0001;
      3'b010: n3582_o = 4'b1100;
      3'b001: n3582_o = 4'b1100;
      default: n3582_o = 4'b1100;
    endcase
  /* decoder.vhd:1569:9  */
  always @*
    case (n3566_o)
      3'b100: n3584_o = 2'b01;
      3'b010: n3584_o = 2'b01;
      3'b001: n3584_o = n3553_o;
      default: n3584_o = 2'b01;
    endcase
  /* decoder.vhd:1568:7  */
  assign n3586_o = opc_mnemonic_s == 6'b101001;
  /* decoder.vhd:1597:13  */
  assign n3588_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1601:13  */
  assign n3593_o = clk_mstate_i == 3'b010;
  assign n3594_o = {n3593_o, n3588_o};
  /* decoder.vhd:1595:11  */
  always @*
    case (n3594_o)
      2'b10: n3597_o = 1'b1;
      2'b01: n3597_o = 1'b0;
      default: n3597_o = 1'b0;
    endcase
  /* decoder.vhd:1595:11  */
  always @*
    case (n3594_o)
      2'b10: n3600_o = 1'b0;
      2'b01: n3600_o = 1'b1;
      default: n3600_o = 1'b0;
    endcase
  /* decoder.vhd:1595:11  */
  always @*
    case (n3594_o)
      2'b10: n3603_o = 1'b1;
      2'b01: n3603_o = 1'b0;
      default: n3603_o = 1'b0;
    endcase
  /* decoder.vhd:1595:11  */
  always @*
    case (n3594_o)
      2'b10: n3606_o = 4'b0001;
      2'b01: n3606_o = 4'b1100;
      default: n3606_o = 4'b1100;
    endcase
  /* decoder.vhd:1594:9  */
  assign n3608_o = clk_second_cycle_i ? n3597_o : 1'b0;
  /* decoder.vhd:1594:9  */
  assign n3610_o = clk_second_cycle_i ? n3600_o : 1'b0;
  /* decoder.vhd:1594:9  */
  assign n3612_o = clk_second_cycle_i ? n3603_o : 1'b0;
  /* decoder.vhd:1594:9  */
  assign n3614_o = clk_second_cycle_i ? n3606_o : 4'b1100;
  /* decoder.vhd:1591:7  */
  assign n3616_o = opc_mnemonic_s == 6'b101010;
  /* decoder.vhd:1615:12  */
  assign n3617_o = ~clk_second_cycle_i;
  /* decoder.vhd:1617:27  */
  assign n3619_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:1618:28  */
  assign n3620_o = opc_opcode_q[1:0];
  /* decoder.vhd:1618:41  */
  assign n3622_o = n3620_o == 2'b00;
  /* decoder.vhd:1620:31  */
  assign n3623_o = opc_opcode_q[1];
  /* decoder.vhd:1620:35  */
  assign n3624_o = ~n3623_o;
  /* decoder.vhd:1620:13  */
  assign n3627_o = n3624_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1620:13  */
  assign n3630_o = n3624_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1620:13  */
  assign n3633_o = n3624_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1620:13  */
  assign n3636_o = n3624_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1618:13  */
  assign n3638_o = n3622_o ? 1'b0 : n3627_o;
  /* decoder.vhd:1618:13  */
  assign n3640_o = n3622_o ? 1'b0 : n3630_o;
  /* decoder.vhd:1618:13  */
  assign n3642_o = n3622_o ? 1'b0 : n3633_o;
  /* decoder.vhd:1618:13  */
  assign n3644_o = n3622_o ? 1'b0 : n3636_o;
  /* decoder.vhd:1618:13  */
  assign n3647_o = n3622_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1617:11  */
  assign n3650_o = n3619_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1617:11  */
  assign n3652_o = n3619_o ? n3638_o : 1'b0;
  /* decoder.vhd:1617:11  */
  assign n3654_o = n3619_o ? n3640_o : 1'b0;
  /* decoder.vhd:1617:11  */
  assign n3656_o = n3619_o ? n3642_o : 1'b0;
  /* decoder.vhd:1617:11  */
  assign n3658_o = n3619_o ? n3644_o : 1'b0;
  /* decoder.vhd:1617:11  */
  assign n3660_o = n3619_o ? n3647_o : 1'b0;
  /* decoder.vhd:1635:13  */
  assign n3662_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1640:13  */
  assign n3664_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1649:30  */
  assign n3665_o = opc_opcode_q[1:0];
  /* decoder.vhd:1649:43  */
  assign n3667_o = n3665_o == 2'b00;
  /* decoder.vhd:1651:33  */
  assign n3668_o = opc_opcode_q[1];
  /* decoder.vhd:1651:37  */
  assign n3669_o = ~n3668_o;
  /* decoder.vhd:1651:15  */
  assign n3672_o = n3669_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1651:15  */
  assign n3675_o = n3669_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1649:15  */
  assign n3678_o = n3667_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1649:15  */
  assign n3680_o = n3667_o ? 1'b0 : n3672_o;
  /* decoder.vhd:1649:15  */
  assign n3682_o = n3667_o ? 1'b0 : n3675_o;
  /* decoder.vhd:1645:13  */
  assign n3684_o = clk_mstate_i == 3'b010;
  assign n3685_o = {n3684_o, n3664_o, n3662_o};
  /* decoder.vhd:1632:11  */
  always @*
    case (n3685_o)
      3'b100: n3689_o = 1'b0;
      3'b010: n3689_o = 1'b1;
      3'b001: n3689_o = 1'b1;
      default: n3689_o = 1'b0;
    endcase
  /* decoder.vhd:1632:11  */
  always @*
    case (n3685_o)
      3'b100: n3693_o = 1'b1;
      3'b010: n3693_o = 1'b1;
      3'b001: n3693_o = 1'b0;
      default: n3693_o = 1'b0;
    endcase
  /* decoder.vhd:1632:11  */
  always @*
    case (n3685_o)
      3'b100: n3695_o = n3678_o;
      3'b010: n3695_o = 1'b0;
      3'b001: n3695_o = 1'b0;
      default: n3695_o = 1'b0;
    endcase
  /* decoder.vhd:1632:11  */
  always @*
    case (n3685_o)
      3'b100: n3697_o = n3680_o;
      3'b010: n3697_o = 1'b0;
      3'b001: n3697_o = 1'b0;
      default: n3697_o = 1'b0;
    endcase
  /* decoder.vhd:1632:11  */
  always @*
    case (n3685_o)
      3'b100: n3699_o = n3682_o;
      3'b010: n3699_o = 1'b0;
      3'b001: n3699_o = 1'b0;
      default: n3699_o = 1'b0;
    endcase
  /* decoder.vhd:1632:11  */
  always @*
    case (n3685_o)
      3'b100: n3702_o = 4'b0001;
      3'b010: n3702_o = 4'b1100;
      3'b001: n3702_o = 4'b1100;
      default: n3702_o = 4'b1100;
    endcase
  /* decoder.vhd:1615:9  */
  assign n3704_o = n3617_o ? 1'b0 : n3689_o;
  /* decoder.vhd:1615:9  */
  assign n3706_o = n3617_o ? n3650_o : 1'b0;
  /* decoder.vhd:1615:9  */
  assign n3708_o = n3617_o ? 1'b0 : n3693_o;
  /* decoder.vhd:1615:9  */
  assign n3710_o = n3617_o ? 1'b0 : n3695_o;
  /* decoder.vhd:1615:9  */
  assign n3712_o = n3617_o ? 1'b0 : n3697_o;
  /* decoder.vhd:1615:9  */
  assign n3714_o = n3617_o ? n3652_o : 1'b0;
  /* decoder.vhd:1615:9  */
  assign n3716_o = n3617_o ? 1'b0 : n3699_o;
  /* decoder.vhd:1615:9  */
  assign n3718_o = n3617_o ? n3654_o : 1'b0;
  /* decoder.vhd:1615:9  */
  assign n3720_o = n3617_o ? 4'b1100 : n3702_o;
  /* decoder.vhd:1615:9  */
  assign n3722_o = n3617_o ? n3656_o : 1'b0;
  /* decoder.vhd:1615:9  */
  assign n3724_o = n3617_o ? n3658_o : 1'b0;
  /* decoder.vhd:1615:9  */
  assign n3726_o = n3617_o ? n3660_o : 1'b0;
  /* decoder.vhd:1612:7  */
  assign n3728_o = opc_mnemonic_s == 6'b101011;
  /* decoder.vhd:1666:24  */
  assign n3729_o = opc_opcode_q[4];
  /* decoder.vhd:1666:28  */
  assign n3730_o = ~n3729_o;
  /* decoder.vhd:1666:9  */
  assign n3733_o = n3730_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1671:12  */
  assign n3734_o = ~clk_second_cycle_i;
  /* decoder.vhd:1671:52  */
  assign n3736_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1671:35  */
  assign n3737_o = n3736_o & n3734_o;
  /* decoder.vhd:1674:26  */
  assign n3738_o = opc_opcode_q[4];
  /* decoder.vhd:1675:28  */
  assign n3739_o = opc_opcode_q[1];
  /* decoder.vhd:1675:32  */
  assign n3740_o = ~n3739_o;
  /* decoder.vhd:1675:13  */
  assign n3743_o = n3740_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1675:13  */
  assign n3746_o = n3740_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1674:11  */
  assign n3749_o = n3738_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1674:11  */
  assign n3751_o = n3738_o ? n3743_o : 1'b0;
  /* decoder.vhd:1674:11  */
  assign n3753_o = n3738_o ? n3746_o : 1'b0;
  /* decoder.vhd:1671:9  */
  assign n3756_o = n3737_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1671:9  */
  assign n3758_o = n3737_o ? n3749_o : 1'b0;
  /* decoder.vhd:1671:9  */
  assign n3760_o = n3737_o ? n3751_o : 1'b0;
  /* decoder.vhd:1671:9  */
  assign n3762_o = n3737_o ? n3753_o : 1'b0;
  /* decoder.vhd:1665:7  */
  assign n3764_o = opc_mnemonic_s == 6'b101101;
  /* decoder.vhd:1690:12  */
  assign n3765_o = ~clk_second_cycle_i;
  /* decoder.vhd:1693:13  */
  assign n3767_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1697:13  */
  assign n3769_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1704:13  */
  assign n3771_o = clk_mstate_i == 3'b100;
  assign n3772_o = {n3771_o, n3769_o, n3767_o};
  /* decoder.vhd:1691:11  */
  always @*
    case (n3772_o)
      3'b100: n3775_o = 1'b1;
      3'b010: n3775_o = 1'b1;
      3'b001: n3775_o = n2073_o;
      default: n3775_o = n2073_o;
    endcase
  /* decoder.vhd:1691:11  */
  always @*
    case (n3772_o)
      3'b100: n3778_o = 1'b1;
      3'b010: n3778_o = 1'b0;
      3'b001: n3778_o = 1'b0;
      default: n3778_o = 1'b0;
    endcase
  /* decoder.vhd:1691:11  */
  always @*
    case (n3772_o)
      3'b100: n3781_o = 1'b1;
      3'b010: n3781_o = 1'b0;
      3'b001: n3781_o = 1'b0;
      default: n3781_o = 1'b0;
    endcase
  /* decoder.vhd:1691:11  */
  always @*
    case (n3772_o)
      3'b100: n3784_o = 1'b0;
      3'b010: n3784_o = 1'b1;
      3'b001: n3784_o = 1'b0;
      default: n3784_o = 1'b0;
    endcase
  /* decoder.vhd:1691:11  */
  always @*
    case (n3772_o)
      3'b100: n3788_o = 2'b11;
      3'b010: n3788_o = 2'b10;
      3'b001: n3788_o = 2'b01;
      default: n3788_o = 2'b01;
    endcase
  /* decoder.vhd:1691:11  */
  always @*
    case (n3772_o)
      3'b100: n3791_o = 1'b0;
      3'b010: n3791_o = 1'b0;
      3'b001: n3791_o = 1'b1;
      default: n3791_o = 1'b0;
    endcase
  /* decoder.vhd:1721:30  */
  assign n3792_o = opc_opcode_q[4];
  /* decoder.vhd:1721:15  */
  assign n3795_o = n3792_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1721:15  */
  assign n3798_o = n3792_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1718:13  */
  assign n3800_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1726:13  */
  assign n3802_o = clk_mstate_i == 3'b001;
  assign n3803_o = {n3802_o, n3800_o};
  /* decoder.vhd:1716:11  */
  always @*
    case (n3803_o)
      2'b10: n3806_o = 1'b0;
      2'b01: n3806_o = 1'b1;
      default: n3806_o = 1'b0;
    endcase
  /* decoder.vhd:1716:11  */
  always @*
    case (n3803_o)
      2'b10: n3809_o = 1'b0;
      2'b01: n3809_o = 1'b1;
      default: n3809_o = 1'b0;
    endcase
  /* decoder.vhd:1716:11  */
  always @*
    case (n3803_o)
      2'b10: n3811_o = 1'b0;
      2'b01: n3811_o = n3795_o;
      default: n3811_o = 1'b0;
    endcase
  /* decoder.vhd:1716:11  */
  always @*
    case (n3803_o)
      2'b10: n3814_o = 1'b1;
      2'b01: n3814_o = 1'b0;
      default: n3814_o = 1'b0;
    endcase
  /* decoder.vhd:1716:11  */
  always @*
    case (n3803_o)
      2'b10: n3816_o = 1'b0;
      2'b01: n3816_o = n3798_o;
      default: n3816_o = 1'b0;
    endcase
  /* decoder.vhd:1690:9  */
  assign n3817_o = n3765_o ? n3775_o : n2073_o;
  /* decoder.vhd:1690:9  */
  assign n3818_o = n3765_o ? n3778_o : n3806_o;
  /* decoder.vhd:1690:9  */
  assign n3820_o = n3765_o ? n3781_o : 1'b0;
  /* decoder.vhd:1690:9  */
  assign n3822_o = n3765_o ? 1'b0 : n3809_o;
  /* decoder.vhd:1690:9  */
  assign n3824_o = n3765_o ? n3784_o : 1'b0;
  /* decoder.vhd:1690:9  */
  assign n3826_o = n3765_o ? 1'b0 : n3811_o;
  /* decoder.vhd:1690:9  */
  assign n3828_o = n3765_o ? n3788_o : 2'b01;
  /* decoder.vhd:1690:9  */
  assign n3830_o = n3765_o ? n3791_o : 1'b0;
  /* decoder.vhd:1690:9  */
  assign n3832_o = n3765_o ? 1'b0 : n3814_o;
  /* decoder.vhd:1690:9  */
  assign n3834_o = n3765_o ? 1'b0 : n3816_o;
  /* decoder.vhd:1689:7  */
  assign n3836_o = opc_mnemonic_s == 6'b101110;
  /* decoder.vhd:1738:25  */
  assign n3838_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1743:26  */
  assign n3839_o = opc_opcode_q[4];
  /* decoder.vhd:1743:11  */
  assign n3842_o = n3839_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1743:11  */
  assign n3844_o = n3839_o ? alu_carry_i : 1'b0;
  /* decoder.vhd:1743:11  */
  assign n3847_o = n3839_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1738:9  */
  assign n3850_o = n3838_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1738:9  */
  assign n3853_o = n3838_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1738:9  */
  assign n3856_o = n3838_o ? 4'b0101 : 4'b1100;
  /* decoder.vhd:1738:9  */
  assign n3858_o = n3838_o ? n3842_o : 1'b0;
  /* decoder.vhd:1738:9  */
  assign n3860_o = n3838_o ? n3844_o : 1'b0;
  /* decoder.vhd:1738:9  */
  assign n3862_o = n3838_o ? n3847_o : 1'b0;
  /* decoder.vhd:1737:7  */
  assign n3864_o = opc_mnemonic_s == 6'b101111;
  /* decoder.vhd:1752:25  */
  assign n3866_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1757:26  */
  assign n3867_o = opc_opcode_q[4];
  /* decoder.vhd:1757:30  */
  assign n3868_o = ~n3867_o;
  /* decoder.vhd:1757:11  */
  assign n3871_o = n3868_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1757:11  */
  assign n3873_o = n3868_o ? alu_carry_i : 1'b0;
  /* decoder.vhd:1757:11  */
  assign n3876_o = n3868_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1752:9  */
  assign n3879_o = n3866_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1752:9  */
  assign n3882_o = n3866_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1752:9  */
  assign n3885_o = n3866_o ? 4'b0110 : 4'b1100;
  /* decoder.vhd:1752:9  */
  assign n3887_o = n3866_o ? n3871_o : 1'b0;
  /* decoder.vhd:1752:9  */
  assign n3889_o = n3866_o ? n3873_o : 1'b0;
  /* decoder.vhd:1752:9  */
  assign n3891_o = n3866_o ? n3876_o : 1'b0;
  /* decoder.vhd:1751:7  */
  assign n3893_o = opc_mnemonic_s == 6'b110000;
  /* decoder.vhd:1766:25  */
  assign n3895_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1767:26  */
  assign n3896_o = opc_opcode_q[4];
  /* decoder.vhd:1767:11  */
  assign n3899_o = n3896_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1767:11  */
  assign n3902_o = n3896_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1766:9  */
  assign n3904_o = n3895_o ? n3899_o : 1'b0;
  /* decoder.vhd:1766:9  */
  assign n3906_o = n3895_o ? n3902_o : 1'b0;
  /* decoder.vhd:1765:7  */
  assign n3908_o = opc_mnemonic_s == 6'b110001;
  /* decoder.vhd:1776:25  */
  assign n3910_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1777:45  */
  assign n3911_o = opc_opcode_q[4];
  /* decoder.vhd:1776:9  */
  assign n3913_o = n3910_o ? n3911_o : 1'b0;
  /* decoder.vhd:1776:9  */
  assign n3916_o = n3910_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1775:7  */
  assign n3918_o = opc_mnemonic_s == 6'b110010;
  /* decoder.vhd:1783:25  */
  assign n3920_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1783:9  */
  assign n3923_o = n3920_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1782:7  */
  assign n3925_o = opc_mnemonic_s == 6'b110011;
  /* decoder.vhd:1789:25  */
  assign n3927_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1790:26  */
  assign n3928_o = opc_opcode_q[4];
  /* decoder.vhd:1790:11  */
  assign n3931_o = n3928_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1790:11  */
  assign n3934_o = n3928_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1789:9  */
  assign n3936_o = n3927_o ? n3931_o : 1'b0;
  /* decoder.vhd:1789:9  */
  assign n3938_o = n3927_o ? n3934_o : 1'b0;
  /* decoder.vhd:1788:7  */
  assign n3940_o = opc_mnemonic_s == 6'b110100;
  /* decoder.vhd:1801:25  */
  assign n3942_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1801:9  */
  assign n3945_o = n3942_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1801:9  */
  assign n3948_o = n3942_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1798:7  */
  assign n3950_o = opc_mnemonic_s == 6'b110101;
  /* decoder.vhd:1812:28  */
  assign n3951_o = opc_opcode_q[3];
  /* decoder.vhd:1812:32  */
  assign n3952_o = ~n3951_o;
  /* decoder.vhd:1811:44  */
  assign n3954_o = 1'b0 | n3952_o;
  /* decoder.vhd:1811:13  */
  assign n3961_o = n3954_o ? 1'b1 : n2073_o;
  /* decoder.vhd:1811:13  */
  assign n3964_o = n3954_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1811:13  */
  assign n3967_o = n3954_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1810:11  */
  assign n3969_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1822:28  */
  assign n3970_o = opc_opcode_q[4];
  /* decoder.vhd:1822:13  */
  assign n3973_o = n3970_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1818:11  */
  assign n3975_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1832:28  */
  assign n3976_o = opc_opcode_q[4];
  /* decoder.vhd:1832:13  */
  assign n3979_o = n3976_o ? 4'b1011 : 4'b1100;
  /* decoder.vhd:1829:11  */
  assign n3981_o = clk_mstate_i == 3'b100;
  assign n3982_o = {n3981_o, n3975_o, n3969_o};
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n3985_o = 1'b0;
      3'b010: n3985_o = 1'b1;
      3'b001: n3985_o = 1'b0;
      default: n3985_o = 1'b0;
    endcase
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n3988_o = 1'b0;
      3'b010: n3988_o = 1'b1;
      3'b001: n3988_o = 1'b0;
      default: n3988_o = 1'b0;
    endcase
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n3991_o = 1'b1;
      3'b010: n3991_o = 1'b0;
      3'b001: n3991_o = 1'b0;
      default: n3991_o = 1'b0;
    endcase
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n3992_o = n2073_o;
      3'b010: n3992_o = n2073_o;
      3'b001: n3992_o = n3961_o;
      default: n3992_o = n2073_o;
    endcase
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n3995_o = 1'b0;
      3'b010: n3995_o = 1'b1;
      3'b001: n3995_o = n3964_o;
      default: n3995_o = 1'b0;
    endcase
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n3997_o = n3979_o;
      3'b010: n3997_o = 4'b1100;
      3'b001: n3997_o = 4'b1100;
      default: n3997_o = 4'b1100;
    endcase
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n3999_o = 1'b0;
      3'b010: n3999_o = n3973_o;
      3'b001: n3999_o = 1'b0;
      default: n3999_o = 1'b0;
    endcase
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n4001_o = 2'b01;
      3'b010: n4001_o = 2'b01;
      3'b001: n4001_o = n3967_o;
      default: n4001_o = 2'b01;
    endcase
  /* decoder.vhd:1808:9  */
  always @*
    case (n3982_o)
      3'b100: n4004_o = 1'b1;
      3'b010: n4004_o = 1'b0;
      3'b001: n4004_o = 1'b0;
      default: n4004_o = 1'b0;
    endcase
  /* decoder.vhd:1807:7  */
  assign n4006_o = opc_mnemonic_s == 6'b110110;
  /* decoder.vhd:1849:28  */
  assign n4007_o = opc_opcode_q[3];
  /* decoder.vhd:1849:32  */
  assign n4008_o = ~n4007_o;
  /* decoder.vhd:1848:44  */
  assign n4010_o = 1'b0 | n4008_o;
  /* decoder.vhd:1848:13  */
  assign n4017_o = n4010_o ? 1'b1 : n2073_o;
  /* decoder.vhd:1848:13  */
  assign n4020_o = n4010_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1848:13  */
  assign n4023_o = n4010_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1847:11  */
  assign n4025_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1854:11  */
  assign n4030_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1858:11  */
  assign n4035_o = clk_mstate_i == 3'b100;
  assign n4036_o = {n4035_o, n4030_o, n4025_o};
  /* decoder.vhd:1845:9  */
  always @*
    case (n4036_o)
      3'b100: n4039_o = 1'b1;
      3'b010: n4039_o = 1'b0;
      3'b001: n4039_o = 1'b0;
      default: n4039_o = 1'b0;
    endcase
  /* decoder.vhd:1845:9  */
  always @*
    case (n4036_o)
      3'b100: n4042_o = 1'b0;
      3'b010: n4042_o = 1'b1;
      3'b001: n4042_o = 1'b0;
      default: n4042_o = 1'b0;
    endcase
  /* decoder.vhd:1845:9  */
  always @*
    case (n4036_o)
      3'b100: n4045_o = 1'b1;
      3'b010: n4045_o = 1'b0;
      3'b001: n4045_o = 1'b0;
      default: n4045_o = 1'b0;
    endcase
  /* decoder.vhd:1845:9  */
  always @*
    case (n4036_o)
      3'b100: n4046_o = n2073_o;
      3'b010: n4046_o = n2073_o;
      3'b001: n4046_o = n4017_o;
      default: n4046_o = n2073_o;
    endcase
  /* decoder.vhd:1845:9  */
  always @*
    case (n4036_o)
      3'b100: n4049_o = 1'b0;
      3'b010: n4049_o = 1'b1;
      3'b001: n4049_o = n4020_o;
      default: n4049_o = 1'b0;
    endcase
  /* decoder.vhd:1845:9  */
  always @*
    case (n4036_o)
      3'b100: n4052_o = 4'b0010;
      3'b010: n4052_o = 4'b1100;
      3'b001: n4052_o = 4'b1100;
      default: n4052_o = 4'b1100;
    endcase
  /* decoder.vhd:1845:9  */
  always @*
    case (n4036_o)
      3'b100: n4054_o = 2'b01;
      3'b010: n4054_o = 2'b01;
      3'b001: n4054_o = n4023_o;
      default: n4054_o = 2'b01;
    endcase
  /* decoder.vhd:1844:7  */
  assign n4056_o = opc_mnemonic_s == 6'b110111;
  /* decoder.vhd:1873:13  */
  assign n4058_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1877:13  */
  assign n4063_o = clk_mstate_i == 3'b010;
  assign n4064_o = {n4063_o, n4058_o};
  /* decoder.vhd:1871:11  */
  always @*
    case (n4064_o)
      2'b10: n4067_o = 1'b1;
      2'b01: n4067_o = 1'b0;
      default: n4067_o = 1'b0;
    endcase
  /* decoder.vhd:1871:11  */
  always @*
    case (n4064_o)
      2'b10: n4070_o = 1'b0;
      2'b01: n4070_o = 1'b1;
      default: n4070_o = 1'b0;
    endcase
  /* decoder.vhd:1871:11  */
  always @*
    case (n4064_o)
      2'b10: n4073_o = 1'b1;
      2'b01: n4073_o = 1'b0;
      default: n4073_o = 1'b0;
    endcase
  /* decoder.vhd:1871:11  */
  always @*
    case (n4064_o)
      2'b10: n4076_o = 4'b0010;
      2'b01: n4076_o = 4'b1100;
      default: n4076_o = 4'b1100;
    endcase
  /* decoder.vhd:1870:9  */
  assign n4078_o = clk_second_cycle_i ? n4067_o : 1'b0;
  /* decoder.vhd:1870:9  */
  assign n4080_o = clk_second_cycle_i ? n4070_o : 1'b0;
  /* decoder.vhd:1870:9  */
  assign n4082_o = clk_second_cycle_i ? n4073_o : 1'b0;
  /* decoder.vhd:1870:9  */
  assign n4084_o = clk_second_cycle_i ? n4076_o : 4'b1100;
  /* decoder.vhd:1867:7  */
  assign n4086_o = opc_mnemonic_s == 6'b111000;
  assign n4087_o = {n4086_o, n4056_o, n4006_o, n3950_o, n3940_o, n3925_o, n3918_o, n3908_o, n3893_o, n3864_o, n3836_o, n3764_o, n3728_o, n3616_o, n3586_o, n3536_o, n3534_o, n3468_o, n3437_o, n3372_o, n3304_o, n3279_o, n3245_o, n3210_o, n3197_o, n3184_o, n3145_o, n3137_o, n3101_o, n3070_o, n3034_o, n3008_o, n2981_o, n2950_o, n2916_o, n2885_o, n2854_o, n2793_o, n2782_o, n2762_o, n2755_o, n2691_o, n2676_o, n2661_o, n2625_o, n2579_o, n2558_o, n2548_o, n2535_o, n2519_o, n2512_o, n2499_o, n2390_o, n2278_o, n2248_o, n2198_o, n2146_o};
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4089_o = n4078_o;
      57'b010000000000000000000000000000000000000000000000000000000: n4089_o = n4039_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4089_o = n3985_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4089_o = n3945_o;
      57'b000010000000000000000000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4089_o = n3879_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4089_o = n3850_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4089_o = n3608_o;
      57'b000000000000001000000000000000000000000000000000000000000: n4089_o = n3569_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4089_o = n3523_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4089_o = n3460_o;
      57'b000000000000000000100000000000000000000000000000000000000: n4089_o = n3425_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4089_o = n3296_o;
      57'b000000000000000000000100000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4089_o = n3189_o;
      57'b000000000000000000000000010000000000000000000000000000000: n4089_o = n3173_o;
      57'b000000000000000000000000001000000000000000000000000000000: n4089_o = n3143_o;
      57'b000000000000000000000000000100000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4089_o = n2837_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4089_o = n2788_o;
      57'b000000000000000000000000000000000000001000000000000000000: n4089_o = n2776_o;
      57'b000000000000000000000000000000000000000100000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4089_o = n2647_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4089_o = n2601_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4089_o = n2540_o;
      57'b000000000000000000000000000000000000000000000000100000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4089_o = n2504_o;
      57'b000000000000000000000000000000000000000000000000000100000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4089_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4089_o = n2270_o;
      57'b000000000000000000000000000000000000000000000000000000100: n4089_o = n2231_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4089_o = n2182_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4089_o = n2119_o;
      default: n4089_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4092_o = n3704_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4092_o = n2839_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4092_o = n2735_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4092_o = n2649_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4092_o = n2603_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4092_o = n2366_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4092_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4092_o = 1'b0;
      default: n4092_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4095_o = n4080_o;
      57'b010000000000000000000000000000000000000000000000000000000: n4095_o = n4042_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4095_o = n3988_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4095_o = n3706_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4095_o = n3610_o;
      57'b000000000000001000000000000000000000000000000000000000000: n4095_o = n3572_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4095_o = n3176_o;
      57'b000000000000000000000000001000000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4095_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4095_o = n2368_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4095_o = n2272_o;
      57'b000000000000000000000000000000000000000000000000000000100: n4095_o = n2234_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4095_o = n2184_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4095_o = n2122_o;
      default: n4095_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4098_o = n4082_o;
      57'b010000000000000000000000000000000000000000000000000000000: n4098_o = n4045_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4098_o = n3991_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4098_o = n3948_o;
      57'b000010000000000000000000000000000000000000000000000000000: n4098_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4098_o = n3882_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4098_o = n3853_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4098_o = n3756_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4098_o = n3708_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4098_o = n3612_o;
      57'b000000000000001000000000000000000000000000000000000000000: n4098_o = n3575_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4098_o = n3524_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4098_o = n3462_o;
      57'b000000000000000000100000000000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4098_o = n3364_o;
      57'b000000000000000000001000000000000000000000000000000000000: n4098_o = n3298_o;
      57'b000000000000000000000100000000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4098_o = n3235_o;
      57'b000000000000000000000001000000000000000000000000000000000: n4098_o = n3202_o;
      57'b000000000000000000000000100000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4098_o = n3127_o;
      57'b000000000000000000000000000010000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4098_o = n3000_o;
      57'b000000000000000000000000000000001000000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4098_o = n2877_o;
      57'b000000000000000000000000000000000000100000000000000000000: n4098_o = n2842_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4098_o = n2737_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4098_o = n2652_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4098_o = n2606_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4098_o = n2543_o;
      57'b000000000000000000000000000000000000000000000000100000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4098_o = n2507_o;
      57'b000000000000000000000000000000000000000000000000000100000: n4098_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4098_o = n2370_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4098_o = n2274_o;
      57'b000000000000000000000000000000000000000000000000000000100: n4098_o = n2237_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4098_o = n2186_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4098_o = n2125_o;
      default: n4098_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4101_o = n3758_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4101_o = n3710_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4101_o = n3525_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4101_o = n2372_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4101_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4101_o = 1'b0;
      default: n4101_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b010000000000000000000000000000000000000000000000000000000: n4103_o = n4046_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4103_o = n3992_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000010000000000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000001000000000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000100000000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000010000000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000001000000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4103_o = n3817_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000001000000000000000000000000000000000000000000: n4103_o = n3576_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000010000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000100000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000001000000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000100000000000000000000000000000000000: n4103_o = n3260_o;
      57'b000000000000000000000010000000000000000000000000000000000: n4103_o = n3236_o;
      57'b000000000000000000000001000000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000100000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000010000000000000000000000000000000: n4103_o = n3177_o;
      57'b000000000000000000000000001000000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000100000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000010000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000001000000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000100000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000010000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000001000000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000100000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000010000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000001000000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000100000000000000000000: n4103_o = n2843_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000001000000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000100000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000010000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000100000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000010000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000010000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000001000000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000000100000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000000010000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000000001000000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000000000100000: n4103_o = n2471_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000000000000100: n4103_o = n2238_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4103_o = n2073_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4103_o = n2126_o;
      default: n4103_o = n2073_o;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4105_o = n4049_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4105_o = n3995_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4105_o = n3818_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4105_o = n3579_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4105_o = n3527_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4105_o = n3269_o;
      57'b000000000000000000000010000000000000000000000000000000000: n4105_o = n3238_o;
      57'b000000000000000000000001000000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4105_o = n3180_o;
      57'b000000000000000000000000001000000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4105_o = n2845_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4105_o = n2739_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4105_o = n2654_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4105_o = n2241_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4105_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4105_o = n2129_o;
      default: n4105_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4108_o = n3760_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4108_o = n3712_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4108_o = n2374_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4108_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4108_o = 1'b0;
      default: n4108_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4111_o = n3714_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4111_o = n2778_o;
      57'b000000000000000000000000000000000000000100000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4111_o = n2376_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4111_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4111_o = 1'b0;
      default: n4111_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4114_o = n3762_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4114_o = n3716_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4114_o = n2378_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4114_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4114_o = 1'b0;
      default: n4114_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4117_o = n3427_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4117_o = n3366_o;
      57'b000000000000000000001000000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4117_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4117_o = 1'b0;
      default: n4117_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4120_o = n3718_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4120_o = n3429_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4120_o = n2780_o;
      57'b000000000000000000000000000000000000000100000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4120_o = n2380_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4120_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4120_o = 1'b0;
      default: n4120_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4123_o = n3431_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4123_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4123_o = 1'b0;
      default: n4123_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4126_o = n3820_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4126_o = n3129_o;
      57'b000000000000000000000000000010000000000000000000000000000: n4126_o = n3093_o;
      57'b000000000000000000000000000001000000000000000000000000000: n4126_o = n3062_o;
      57'b000000000000000000000000000000100000000000000000000000000: n4126_o = n3028_o;
      57'b000000000000000000000000000000010000000000000000000000000: n4126_o = n3002_o;
      57'b000000000000000000000000000000001000000000000000000000000: n4126_o = n2973_o;
      57'b000000000000000000000000000000000100000000000000000000000: n4126_o = n2942_o;
      57'b000000000000000000000000000000000010000000000000000000000: n4126_o = n2908_o;
      57'b000000000000000000000000000000000001000000000000000000000: n4126_o = n2879_o;
      57'b000000000000000000000000000000000000100000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4126_o = n2741_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4126_o = n2473_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4126_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4126_o = 1'b0;
      default: n4126_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4129_o = n2475_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4129_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4129_o = 1'b0;
      default: n4129_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4132_o = n3822_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4132_o = n2975_o;
      57'b000000000000000000000000000000000100000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4132_o = n2477_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4132_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4132_o = 1'b0;
      default: n4132_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4135_o = n2479_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4135_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4135_o = 1'b0;
      default: n4135_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4138_o = n3192_o;
      57'b000000000000000000000000010000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4138_o = n2481_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4138_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4138_o = 1'b0;
      default: n4138_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4141_o = n3824_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4141_o = n3195_o;
      57'b000000000000000000000000010000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4141_o = n2483_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4141_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4141_o = 1'b0;
      default: n4141_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4144_o = n3826_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4144_o = n3205_o;
      57'b000000000000000000000000100000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4144_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4144_o = 1'b0;
      default: n4144_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4147_o = n3208_o;
      57'b000000000000000000000000100000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4147_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4147_o = 1'b0;
      default: n4147_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4151_o = n4084_o;
      57'b010000000000000000000000000000000000000000000000000000000: n4151_o = n4052_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4151_o = n3997_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4151_o = 4'b0111;
      57'b000010000000000000000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000001000000000000000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000100000000000000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000010000000000000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000001000000000000000000000000000000000000000000000000: n4151_o = n3885_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4151_o = n3856_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000001000000000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000100000000000000000000000000000000000000000000: n4151_o = n3720_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4151_o = n3614_o;
      57'b000000000000001000000000000000000000000000000000000000000: n4151_o = n3582_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000010000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000001000000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000100000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000010000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000001000000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000100000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000010000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000001000000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000100000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000010000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000001000000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000100000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000010000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000001000000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000100000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000010000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000001000000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000100000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000010000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000001000000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000100000000000000000000: n4151_o = n2848_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000001000000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000100000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000010000000000000000: n4151_o = n2743_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000000100000000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000000010000000000000: n4151_o = n2657_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4151_o = n2608_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000000000010000000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000000000001000000000: n4151_o = n2546_o;
      57'b000000000000000000000000000000000000000000000000100000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000000000000010000000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000000000000001000000: n4151_o = n2510_o;
      57'b000000000000000000000000000000000000000000000000000100000: n4151_o = 4'b1100;
      57'b000000000000000000000000000000000000000000000000000010000: n4151_o = n2382_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4151_o = n2276_o;
      57'b000000000000000000000000000000000000000000000000000000100: n4151_o = n2244_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4151_o = n2188_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4151_o = n2132_o;
      default: n4151_o = 4'b1100;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4154_o = n3887_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4154_o = n3858_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4154_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4154_o = n2190_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4154_o = n2134_o;
      default: n4154_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4157_o = n2612_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4157_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4157_o = 1'b0;
      default: n4157_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4160_o = n3999_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4160_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4160_o = 1'b0;
      default: n4160_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4163_o = n2615_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4163_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4163_o = 1'b0;
      default: n4163_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4166_o = n2618_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4166_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4166_o = 1'b0;
      default: n4166_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4170_o = 1'b1;
      57'b000000000000000001000000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4170_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4170_o = 1'b0;
      default: n4170_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4175_o = 1'b1;
      57'b000000000000000000010000000000000000000000000000000000000: n4175_o = 1'b1;
      57'b000000000000000000001000000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4175_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4175_o = 1'b0;
      default: n4175_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4179_o = n3473_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4179_o = 1'b1;
      57'b000000000000000000000000000000000000001000000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4179_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4179_o = 1'b0;
      default: n4179_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4182_o = n3733_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4182_o = n3476_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4182_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4182_o = 1'b0;
      default: n4182_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4185_o = n3131_o;
      57'b000000000000000000000000000010000000000000000000000000000: n4185_o = n3095_o;
      57'b000000000000000000000000000001000000000000000000000000000: n4185_o = n3064_o;
      57'b000000000000000000000000000000100000000000000000000000000: n4185_o = n3030_o;
      57'b000000000000000000000000000000010000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4185_o = n2944_o;
      57'b000000000000000000000000000000000010000000000000000000000: n4185_o = n2910_o;
      57'b000000000000000000000000000000000001000000000000000000000: n4185_o = n2881_o;
      57'b000000000000000000000000000000000000100000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4185_o = n2745_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4185_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4185_o = 1'b0;
      default: n4185_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b010000000000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b001000000000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000100000000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000010000000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000001000000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000100000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000010000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000001000000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000100000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000010000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000001000000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000100000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000010000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000001000000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000100000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000010000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000001000000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000100000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000010000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000001000000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000100000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000010000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000001000000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000100000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000010000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000001000000000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000100000000000000000000000000000: n4193_o = 4'b0001;
      57'b000000000000000000000000000010000000000000000000000000000: n4193_o = 4'b1000;
      57'b000000000000000000000000000001000000000000000000000000000: n4193_o = n3039_o;
      57'b000000000000000000000000000000100000000000000000000000000: n4193_o = 4'b0101;
      57'b000000000000000000000000000000010000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000001000000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000100000000000000000000000: n4193_o = n2946_o;
      57'b000000000000000000000000000000000010000000000000000000000: n4193_o = 4'b0010;
      57'b000000000000000000000000000000000001000000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000100000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000010000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000001000000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000100000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000010000000000000000: n4193_o = n2747_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000100000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000010000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000001000000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000100000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000010000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000001000000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000100000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000010000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000001000000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000000100000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000000010000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000000001000: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000000000100: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000000000010: n4193_o = 4'b0000;
      57'b000000000000000000000000000000000000000000000000000000001: n4193_o = 4'b0000;
      default: n4193_o = 4'b0000;
    endcase
  assign n4195_o = opc_opcode_q[5];
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b010000000000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000010000000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000001000000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000100000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000010000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000001000000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000001000000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000010000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000100000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000001000000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000100000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000010000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000001000000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000100000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000010000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000001000000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000100000000000000000000000000000: n4196_o = n3113_o;
      57'b000000000000000000000000000010000000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000001000000000000000000000000000: n4196_o = n3048_o;
      57'b000000000000000000000000000000100000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000010000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000001000000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000100000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000010000000000000000000000: n4196_o = n2894_o;
      57'b000000000000000000000000000000000001000000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000100000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000001000000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000100000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000010000000000000000: n4196_o = n2749_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000100000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000010000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000010000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000001000000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000100000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000010000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000001000000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000000100000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000000000100: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4196_o = n4195_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4196_o = n4195_o;
      default: n4196_o = n4195_o;
    endcase
  assign n4197_o = opc_opcode_q[7:6];
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b010000000000000000000000000000000000000000000000000000000: n4199_o = n4054_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4199_o = n4001_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000010000000000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000001000000000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000100000000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000010000000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000001000000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000100000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000010000000000000000000000000000000000000000000000: n4199_o = n3828_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000100000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000010000000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000001000000000000000000000000000000000000000000: n4199_o = n3584_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000010000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000001000000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000100000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000010000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000001000000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000100000000000000000000000000000000000: n4199_o = n3271_o;
      57'b000000000000000000000010000000000000000000000000000000000: n4199_o = n3240_o;
      57'b000000000000000000000001000000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000100000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000010000000000000000000000000000000: n4199_o = n3182_o;
      57'b000000000000000000000000001000000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000100000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000010000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000001000000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000100000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000010000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000001000000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000100000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000010000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000001000000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000100000000000000000000: n4199_o = n2850_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000001000000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000100000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000010000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000001000000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000100000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000010000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000001000000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000100000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000010000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000001000000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000000100000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000000010000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000000001000000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000000000100000: n4199_o = n2485_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000000000001000: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000000000000100: n4199_o = n2246_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4199_o = 2'b01;
      57'b000000000000000000000000000000000000000000000000000000001: n4199_o = n2136_o;
      default: n4199_o = 2'b01;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4202_o = n3722_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4202_o = n2384_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4202_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4202_o = 1'b0;
      default: n4202_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4205_o = n3724_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4205_o = n2386_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4205_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4205_o = 1'b0;
      default: n4205_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b010000000000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b001000000000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000100000000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000010000000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000001000000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000100000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000010000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000001000000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000100000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000010000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000001000000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000100000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000010000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000001000000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000100000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000010000000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000001000000000000000000000000000000000000000: n4208_o = n3464_o;
      57'b000000000000000000100000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000010000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000001000000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000100000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000010000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000001000000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000100000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000010000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000001000000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000100000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000010000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000001000000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000100000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000010000000000000000000000000: n4208_o = n3004_o;
      57'b000000000000000000000000000000001000000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000100000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000010000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000001000000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000100000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000010000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000001000000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000100000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000010000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000001000000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000100000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000010000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000001000000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000100000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000010000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000001000000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000100000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000010000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000001000000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000000100000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000000010000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000000001000: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000000000100: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000000000010: n4208_o = 2'b00;
      57'b000000000000000000000000000000000000000000000000000000001: n4208_o = 2'b00;
      default: n4208_o = 2'b00;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4211_o = n3913_o;
      57'b000000010000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4211_o = n3889_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4211_o = n3860_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4211_o = n2620_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4211_o = n2573_o;
      57'b000000000000000000000000000000000000000000000010000000000: n4211_o = n2553_o;
      57'b000000000000000000000000000000000000000000000001000000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4211_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4211_o = n2192_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4211_o = n2138_o;
      default: n4211_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4214_o = n2487_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4214_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4214_o = 1'b0;
      default: n4214_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4217_o = n3830_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4217_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4217_o = 1'b0;
      default: n4217_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4220_o = n3891_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4220_o = n3862_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4220_o = n2623_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4220_o = n2556_o;
      57'b000000000000000000000000000000000000000000000001000000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4220_o = n2517_o;
      57'b000000000000000000000000000000000000000000000000001000000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4220_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4220_o = n2194_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4220_o = n2141_o;
      default: n4220_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4223_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4223_o = n2196_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4223_o = n2144_o;
      default: n4223_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4226_o = n2575_o;
      57'b000000000000000000000000000000000000000000000010000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4226_o = n2531_o;
      57'b000000000000000000000000000000000000000000000000010000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4226_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4226_o = 1'b0;
      default: n4226_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4229_o = n3916_o;
      57'b000000010000000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4229_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4229_o = 1'b0;
      default: n4229_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4232_o = n3300_o;
      57'b000000000000000000000100000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4232_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4232_o = 1'b0;
      default: n4232_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4235_o = n3302_o;
      57'b000000000000000000000100000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4235_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4235_o = 1'b0;
      default: n4235_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4238_o = n3936_o;
      57'b000001000000000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4238_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4238_o = 1'b0;
      default: n4238_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4241_o = n3938_o;
      57'b000001000000000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4241_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4241_o = 1'b0;
      default: n4241_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4244_o = n3923_o;
      57'b000000100000000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4244_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4244_o = 1'b0;
      default: n4244_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4267_o = 1'b1;
      57'b010000000000000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000010000000000000000000000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000001000000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000100000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000010000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000100000000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000010000000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000001000000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000000100000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000000010000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000000001000000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000000000100000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000000000010000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000000000001000000000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000000000000100000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4267_o = 1'b1;
      57'b000000000000000000000000000000000000000001000000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4267_o = 1'b1;
      57'b000000000000000000000000000000000000000000000000000010000: n4267_o = 1'b1;
      57'b000000000000000000000000000000000000000000000000000001000: n4267_o = 1'b1;
      57'b000000000000000000000000000000000000000000000000000000100: n4267_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4267_o = 1'b1;
      57'b000000000000000000000000000000000000000000000000000000001: n4267_o = 1'b0;
      default: n4267_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4270_o = n3466_o;
      57'b000000000000000000100000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4270_o = n3135_o;
      57'b000000000000000000000000000010000000000000000000000000000: n4270_o = n3097_o;
      57'b000000000000000000000000000001000000000000000000000000000: n4270_o = n3068_o;
      57'b000000000000000000000000000000100000000000000000000000000: n4270_o = n3032_o;
      57'b000000000000000000000000000000010000000000000000000000000: n4270_o = n3006_o;
      57'b000000000000000000000000000000001000000000000000000000000: n4270_o = n2977_o;
      57'b000000000000000000000000000000000100000000000000000000000: n4270_o = n2948_o;
      57'b000000000000000000000000000000000010000000000000000000000: n4270_o = n2914_o;
      57'b000000000000000000000000000000000001000000000000000000000: n4270_o = n2883_o;
      57'b000000000000000000000000000000000000100000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4270_o = n2751_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4270_o = n2489_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4270_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4270_o = 1'b0;
      default: n4270_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4273_o = n2491_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4273_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4273_o = 1'b0;
      default: n4273_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4276_o = n3832_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4276_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4276_o = 1'b0;
      default: n4276_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4279_o = n2533_o;
      57'b000000000000000000000000000000000000000000000000010000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4279_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4279_o = 1'b0;
      default: n4279_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4282_o = n2577_o;
      57'b000000000000000000000000000000000000000000000010000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4282_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4282_o = 1'b0;
      default: n4282_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4285_o = n3904_o;
      57'b000000001000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4285_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4285_o = 1'b0;
      default: n4285_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4288_o = n3906_o;
      57'b000000001000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4288_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4288_o = 1'b0;
      default: n4288_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4291_o = n2760_o;
      57'b000000000000000000000000000000000000000010000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4291_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4291_o = 1'b0;
      default: n4291_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b010000000000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000010000000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000001000000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000100000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000010000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000001000000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000001000000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000010000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000100000000000000000000000000000000000000: n4293_o = n3433_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4293_o = n3368_o;
      57'b000000000000000000001000000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000100000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000010000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000001000000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000100000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000010000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000001000000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000100000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000010000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000001000000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000100000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000010000000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000001000000000000000000000000: n4293_o = n2978_o;
      57'b000000000000000000000000000000000100000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000010000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000001000000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000100000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000001000000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000100000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000010000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000100000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000010000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000010000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000001000000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000000100000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000000010000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000000001000000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000000000100000: n4293_o = n2492_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000000000000100: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4293_o = n2077_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4293_o = n2077_o;
      default: n4293_o = n2077_o;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b010000000000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b001000000000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000010000000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000001000000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000100000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000010000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000001000000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000100000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000010000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000100000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000001000000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000100000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000010000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000100000000000000000000000000000000000000: n4294_o = n3434_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4294_o = n3369_o;
      57'b000000000000000000001000000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000100000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000010000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000001000000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000100000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000010000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000001000000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000100000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000010000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000001000000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000100000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000010000000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000001000000000000000000000000: n4294_o = n2979_o;
      57'b000000000000000000000000000000000100000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000010000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000001000000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000100000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000001000000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000100000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000010000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000100000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000010000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000100000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000010000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000001000000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000000100000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000000010000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000000001000000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000000000100000: n4294_o = n2493_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000000000000100: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000000000000010: n4294_o = n2081_o;
      57'b000000000000000000000000000000000000000000000000000000001: n4294_o = n2081_o;
      default: n4294_o = n2081_o;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4296_o = n3726_o;
      57'b000000000000010000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4296_o = n3529_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4296_o = n2791_o;
      57'b000000000000000000000000000000000000001000000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4296_o = n2388_o;
      57'b000000000000000000000000000000000000000000000000000001000: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4296_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4296_o = 1'b0;
      default: n4296_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4299_o = n4004_o;
      57'b000100000000000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4299_o = n3277_o;
      57'b000000000000000000000010000000000000000000000000000000000: n4299_o = n3243_o;
      57'b000000000000000000000001000000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4299_o = n2852_o;
      57'b000000000000000000000000000000000000010000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4299_o = n2753_o;
      57'b000000000000000000000000000000000000000001000000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4299_o = n2659_o;
      57'b000000000000000000000000000000000000000000001000000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4299_o = n2495_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4299_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4299_o = 1'b0;
      default: n4299_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4302_o = n3435_o;
      57'b000000000000000000010000000000000000000000000000000000000: n4302_o = n3370_o;
      57'b000000000000000000001000000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4302_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4302_o = 1'b0;
      default: n4302_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4305_o = n3532_o;
      57'b000000000000000001000000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4305_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4305_o = 1'b0;
      default: n4305_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4308_o = n3099_o;
      57'b000000000000000000000000000001000000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4308_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4308_o = 1'b0;
      default: n4308_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4311_o = n2687_o;
      57'b000000000000000000000000000000000000000000100000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4311_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4311_o = 1'b0;
      default: n4311_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4314_o = n2689_o;
      57'b000000000000000000000000000000000000000000100000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4314_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4314_o = 1'b0;
      default: n4314_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4317_o = n2672_o;
      57'b000000000000000000000000000000000000000000010000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4317_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4317_o = 1'b0;
      default: n4317_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4320_o = n2674_o;
      57'b000000000000000000000000000000000000000000010000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4320_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4320_o = 1'b0;
      default: n4320_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4323_o = n3834_o;
      57'b000000000001000000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000010000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4323_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4323_o = 1'b0;
      default: n4323_o = 1'b0;
    endcase
  /* decoder.vhd:606:5  */
  always @*
    case (n4087_o)
      57'b100000000000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b010000000000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b001000000000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000100000000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000010000000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000001000000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000100000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000010000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000001000000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000100000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000010000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000001000000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000100000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000010000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000001000000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000100000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000010000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000001000000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000100000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000010000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000001000000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000100000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000010000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000001000000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000100000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000010000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000001000000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000100000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000010000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000001000000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000100000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000010000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000001000000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000100000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000010000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000001000000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000100000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000010000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000001000000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000100000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000010000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000001000000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000100000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000010000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000001000000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000100000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000010000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000001000000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000100000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000010000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000001000000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000100000: n4326_o = n2497_o;
      57'b000000000000000000000000000000000000000000000000000010000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000001000: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000100: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000010: n4326_o = 1'b0;
      57'b000000000000000000000000000000000000000000000000000000001: n4326_o = 1'b0;
      default: n4326_o = 1'b0;
    endcase
  /* decoder.vhd:1912:14  */
  assign n4330_o = ~res_i;
  /* decoder.vhd:1929:28  */
  assign n4333_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:1929:9  */
  assign n4335_o = n4333_o ? 1'b0 : branch_taken_q;
  /* decoder.vhd:1927:9  */
  assign n4337_o = branch_taken_s ? 1'b1 : n4335_o;
  /* decoder.vhd:1938:27  */
  assign n4338_o = ~f1_q;
  /* decoder.vhd:1937:9  */
  assign n4339_o = cpl_f1_s ? n4338_o : f1_q;
  /* decoder.vhd:1935:9  */
  assign n4341_o = clear_f1_s ? 1'b0 : n4339_o;
  /* decoder.vhd:1944:9  */
  assign n4343_o = set_mb_s ? 1'b1 : mb_q;
  /* decoder.vhd:1942:9  */
  assign n4345_o = clear_mb_s ? 1'b0 : n4343_o;
  /* decoder.vhd:1924:7  */
  assign n4351_o = en_clk_i & ent0_clk_s;
  /* decoder.vhd:2000:27  */
  assign n4365_o = read_dec_s ? data_s : 8'b11111111;
  /* decoder.vhd:2002:48  */
  assign n4367_o = en_clk_i & dm_write_dmem_s;
  /* decoder.vhd:2003:48  */
  assign n4368_o = pm_inc_pc_s | add_inc_pc_s;
  /* decoder.vhd:2004:48  */
  assign n4369_o = pm_write_pmem_addr_s | add_write_pmem_addr_s;
  /* decoder.vhd:2006:48  */
  assign n4370_o = bus_read_bus_s | add_read_bus_s;
  /* decoder.vhd:280:5  */
  assign n4371_o = en_clk_i ? n1912_o : opc_opcode_q;
  /* decoder.vhd:280:5  */
  always @(posedge clk_i or posedge n1906_o)
    if (n1906_o)
      n4372_q <= 8'b00000000;
    else
      n4372_q <= n4371_o;
  /* decoder.vhd:1923:5  */
  assign n4373_o = en_clk_i ? n4337_o : branch_taken_q;
  /* decoder.vhd:1923:5  */
  always @(posedge clk_i or posedge n4330_o)
    if (n4330_o)
      n4374_q <= 1'b0;
    else
      n4374_q <= n4373_o;
  /* decoder.vhd:1923:5  */
  assign n4375_o = en_clk_i ? n4341_o : f1_q;
  /* decoder.vhd:1923:5  */
  always @(posedge clk_i or posedge n4330_o)
    if (n4330_o)
      n4376_q <= 1'b0;
    else
      n4376_q <= n4375_o;
  /* decoder.vhd:1923:5  */
  assign n4377_o = en_clk_i ? n4345_o : mb_q;
  /* decoder.vhd:1923:5  */
  always @(posedge clk_i or posedge n4330_o)
    if (n4330_o)
      n4378_q <= 1'b0;
    else
      n4378_q <= n4377_o;
  /* decoder.vhd:1923:5  */
  assign n4379_o = n4351_o ? 1'b1 : t0_dir_q;
  /* decoder.vhd:1923:5  */
  always @(posedge clk_i or posedge n4330_o)
    if (n4330_o)
      n4380_q <= 1'b0;
    else
      n4380_q <= n4379_o;
  /* decoder.vhd:280:5  */
  assign n4381_o = en_clk_i ? n1913_o : mnemonic_q;
  /* decoder.vhd:280:5  */
  always @(posedge clk_i or posedge n1906_o)
    if (n1906_o)
      n4382_q <= 6'b101000;
    else
      n4382_q <= n4381_o;
  /* decoder.vhd:276:5  */
  assign n4383_o = {n4197_o, n4196_o};
endmodule